// This is the unpowered netlist.
module audiodac (clk_i,
    ds_n_o,
    ds_o,
    fifo_ack_o,
    fifo_empty_o,
    fifo_full_o,
    fifo_rdy_i,
    mode_i,
    rst_n_i,
    tst_fifo_loop_i,
    tst_sinegen_en_i,
    fifo_i,
    osr_i,
    tst_sinegen_step_i,
    volume_i);
 input clk_i;
 output ds_n_o;
 output ds_o;
 output fifo_ack_o;
 output fifo_empty_o;
 output fifo_full_o;
 input fifo_rdy_i;
 input mode_i;
 input rst_n_i;
 input tst_fifo_loop_i;
 input tst_sinegen_en_i;
 input [15:0] fifo_i;
 input [1:0] osr_i;
 input [5:0] tst_sinegen_step_i;
 input [3:0] volume_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire \dsmod0.accu1[0] ;
 wire \dsmod0.accu1[10] ;
 wire \dsmod0.accu1[11] ;
 wire \dsmod0.accu1[12] ;
 wire \dsmod0.accu1[13] ;
 wire \dsmod0.accu1[14] ;
 wire \dsmod0.accu1[15] ;
 wire \dsmod0.accu1[1] ;
 wire \dsmod0.accu1[2] ;
 wire \dsmod0.accu1[3] ;
 wire \dsmod0.accu1[4] ;
 wire \dsmod0.accu1[5] ;
 wire \dsmod0.accu1[6] ;
 wire \dsmod0.accu1[7] ;
 wire \dsmod0.accu1[8] ;
 wire \dsmod0.accu1[9] ;
 wire \dsmod0.accu2[0] ;
 wire \dsmod0.accu2[10] ;
 wire \dsmod0.accu2[11] ;
 wire \dsmod0.accu2[12] ;
 wire \dsmod0.accu2[13] ;
 wire \dsmod0.accu2[14] ;
 wire \dsmod0.accu2[15] ;
 wire \dsmod0.accu2[1] ;
 wire \dsmod0.accu2[2] ;
 wire \dsmod0.accu2[3] ;
 wire \dsmod0.accu2[4] ;
 wire \dsmod0.accu2[5] ;
 wire \dsmod0.accu2[6] ;
 wire \dsmod0.accu2[7] ;
 wire \dsmod0.accu2[8] ;
 wire \dsmod0.accu2[9] ;
 wire \dsmod0.accu3[0] ;
 wire \dsmod0.accu3[1] ;
 wire \dsmod0.fetch_ctr[0] ;
 wire \dsmod0.fetch_ctr[1] ;
 wire \dsmod0.fetch_ctr[2] ;
 wire \dsmod0.fetch_ctr[3] ;
 wire \dsmod0.fetch_ctr[4] ;
 wire \dsmod0.fetch_ctr[5] ;
 wire \dsmod0.fetch_ctr[6] ;
 wire \dsmod0.fetch_ctr[7] ;
 wire \dsmod0.mod2_ctr[0] ;
 wire \dsmod0.mod2_ctr[1] ;
 wire \dsmod0.mod2_out[0] ;
 wire \dsmod0.mod2_out[1] ;
 wire \fifo0.fifo_data[0] ;
 wire \fifo0.fifo_data[10] ;
 wire \fifo0.fifo_data[11] ;
 wire \fifo0.fifo_data[12] ;
 wire \fifo0.fifo_data[13] ;
 wire \fifo0.fifo_data[14] ;
 wire \fifo0.fifo_data[15] ;
 wire \fifo0.fifo_data[1] ;
 wire \fifo0.fifo_data[2] ;
 wire \fifo0.fifo_data[3] ;
 wire \fifo0.fifo_data[4] ;
 wire \fifo0.fifo_data[5] ;
 wire \fifo0.fifo_data[6] ;
 wire \fifo0.fifo_data[7] ;
 wire \fifo0.fifo_data[8] ;
 wire \fifo0.fifo_data[9] ;
 wire \fifo0.fifo_data_del1[0] ;
 wire \fifo0.fifo_data_del1[10] ;
 wire \fifo0.fifo_data_del1[11] ;
 wire \fifo0.fifo_data_del1[12] ;
 wire \fifo0.fifo_data_del1[13] ;
 wire \fifo0.fifo_data_del1[14] ;
 wire \fifo0.fifo_data_del1[15] ;
 wire \fifo0.fifo_data_del1[1] ;
 wire \fifo0.fifo_data_del1[2] ;
 wire \fifo0.fifo_data_del1[3] ;
 wire \fifo0.fifo_data_del1[4] ;
 wire \fifo0.fifo_data_del1[5] ;
 wire \fifo0.fifo_data_del1[6] ;
 wire \fifo0.fifo_data_del1[7] ;
 wire \fifo0.fifo_data_del1[8] ;
 wire \fifo0.fifo_data_del1[9] ;
 wire \fifo0.fifo_rdy ;
 wire \fifo0.fifo_rdy_del1 ;
 wire \fifo0.fifo_store[0][0] ;
 wire \fifo0.fifo_store[0][10] ;
 wire \fifo0.fifo_store[0][11] ;
 wire \fifo0.fifo_store[0][12] ;
 wire \fifo0.fifo_store[0][13] ;
 wire \fifo0.fifo_store[0][14] ;
 wire \fifo0.fifo_store[0][15] ;
 wire \fifo0.fifo_store[0][1] ;
 wire \fifo0.fifo_store[0][2] ;
 wire \fifo0.fifo_store[0][3] ;
 wire \fifo0.fifo_store[0][4] ;
 wire \fifo0.fifo_store[0][5] ;
 wire \fifo0.fifo_store[0][6] ;
 wire \fifo0.fifo_store[0][7] ;
 wire \fifo0.fifo_store[0][8] ;
 wire \fifo0.fifo_store[0][9] ;
 wire \fifo0.fifo_store[100][0] ;
 wire \fifo0.fifo_store[100][10] ;
 wire \fifo0.fifo_store[100][11] ;
 wire \fifo0.fifo_store[100][12] ;
 wire \fifo0.fifo_store[100][13] ;
 wire \fifo0.fifo_store[100][14] ;
 wire \fifo0.fifo_store[100][15] ;
 wire \fifo0.fifo_store[100][1] ;
 wire \fifo0.fifo_store[100][2] ;
 wire \fifo0.fifo_store[100][3] ;
 wire \fifo0.fifo_store[100][4] ;
 wire \fifo0.fifo_store[100][5] ;
 wire \fifo0.fifo_store[100][6] ;
 wire \fifo0.fifo_store[100][7] ;
 wire \fifo0.fifo_store[100][8] ;
 wire \fifo0.fifo_store[100][9] ;
 wire \fifo0.fifo_store[101][0] ;
 wire \fifo0.fifo_store[101][10] ;
 wire \fifo0.fifo_store[101][11] ;
 wire \fifo0.fifo_store[101][12] ;
 wire \fifo0.fifo_store[101][13] ;
 wire \fifo0.fifo_store[101][14] ;
 wire \fifo0.fifo_store[101][15] ;
 wire \fifo0.fifo_store[101][1] ;
 wire \fifo0.fifo_store[101][2] ;
 wire \fifo0.fifo_store[101][3] ;
 wire \fifo0.fifo_store[101][4] ;
 wire \fifo0.fifo_store[101][5] ;
 wire \fifo0.fifo_store[101][6] ;
 wire \fifo0.fifo_store[101][7] ;
 wire \fifo0.fifo_store[101][8] ;
 wire \fifo0.fifo_store[101][9] ;
 wire \fifo0.fifo_store[102][0] ;
 wire \fifo0.fifo_store[102][10] ;
 wire \fifo0.fifo_store[102][11] ;
 wire \fifo0.fifo_store[102][12] ;
 wire \fifo0.fifo_store[102][13] ;
 wire \fifo0.fifo_store[102][14] ;
 wire \fifo0.fifo_store[102][15] ;
 wire \fifo0.fifo_store[102][1] ;
 wire \fifo0.fifo_store[102][2] ;
 wire \fifo0.fifo_store[102][3] ;
 wire \fifo0.fifo_store[102][4] ;
 wire \fifo0.fifo_store[102][5] ;
 wire \fifo0.fifo_store[102][6] ;
 wire \fifo0.fifo_store[102][7] ;
 wire \fifo0.fifo_store[102][8] ;
 wire \fifo0.fifo_store[102][9] ;
 wire \fifo0.fifo_store[103][0] ;
 wire \fifo0.fifo_store[103][10] ;
 wire \fifo0.fifo_store[103][11] ;
 wire \fifo0.fifo_store[103][12] ;
 wire \fifo0.fifo_store[103][13] ;
 wire \fifo0.fifo_store[103][14] ;
 wire \fifo0.fifo_store[103][15] ;
 wire \fifo0.fifo_store[103][1] ;
 wire \fifo0.fifo_store[103][2] ;
 wire \fifo0.fifo_store[103][3] ;
 wire \fifo0.fifo_store[103][4] ;
 wire \fifo0.fifo_store[103][5] ;
 wire \fifo0.fifo_store[103][6] ;
 wire \fifo0.fifo_store[103][7] ;
 wire \fifo0.fifo_store[103][8] ;
 wire \fifo0.fifo_store[103][9] ;
 wire \fifo0.fifo_store[104][0] ;
 wire \fifo0.fifo_store[104][10] ;
 wire \fifo0.fifo_store[104][11] ;
 wire \fifo0.fifo_store[104][12] ;
 wire \fifo0.fifo_store[104][13] ;
 wire \fifo0.fifo_store[104][14] ;
 wire \fifo0.fifo_store[104][15] ;
 wire \fifo0.fifo_store[104][1] ;
 wire \fifo0.fifo_store[104][2] ;
 wire \fifo0.fifo_store[104][3] ;
 wire \fifo0.fifo_store[104][4] ;
 wire \fifo0.fifo_store[104][5] ;
 wire \fifo0.fifo_store[104][6] ;
 wire \fifo0.fifo_store[104][7] ;
 wire \fifo0.fifo_store[104][8] ;
 wire \fifo0.fifo_store[104][9] ;
 wire \fifo0.fifo_store[105][0] ;
 wire \fifo0.fifo_store[105][10] ;
 wire \fifo0.fifo_store[105][11] ;
 wire \fifo0.fifo_store[105][12] ;
 wire \fifo0.fifo_store[105][13] ;
 wire \fifo0.fifo_store[105][14] ;
 wire \fifo0.fifo_store[105][15] ;
 wire \fifo0.fifo_store[105][1] ;
 wire \fifo0.fifo_store[105][2] ;
 wire \fifo0.fifo_store[105][3] ;
 wire \fifo0.fifo_store[105][4] ;
 wire \fifo0.fifo_store[105][5] ;
 wire \fifo0.fifo_store[105][6] ;
 wire \fifo0.fifo_store[105][7] ;
 wire \fifo0.fifo_store[105][8] ;
 wire \fifo0.fifo_store[105][9] ;
 wire \fifo0.fifo_store[106][0] ;
 wire \fifo0.fifo_store[106][10] ;
 wire \fifo0.fifo_store[106][11] ;
 wire \fifo0.fifo_store[106][12] ;
 wire \fifo0.fifo_store[106][13] ;
 wire \fifo0.fifo_store[106][14] ;
 wire \fifo0.fifo_store[106][15] ;
 wire \fifo0.fifo_store[106][1] ;
 wire \fifo0.fifo_store[106][2] ;
 wire \fifo0.fifo_store[106][3] ;
 wire \fifo0.fifo_store[106][4] ;
 wire \fifo0.fifo_store[106][5] ;
 wire \fifo0.fifo_store[106][6] ;
 wire \fifo0.fifo_store[106][7] ;
 wire \fifo0.fifo_store[106][8] ;
 wire \fifo0.fifo_store[106][9] ;
 wire \fifo0.fifo_store[107][0] ;
 wire \fifo0.fifo_store[107][10] ;
 wire \fifo0.fifo_store[107][11] ;
 wire \fifo0.fifo_store[107][12] ;
 wire \fifo0.fifo_store[107][13] ;
 wire \fifo0.fifo_store[107][14] ;
 wire \fifo0.fifo_store[107][15] ;
 wire \fifo0.fifo_store[107][1] ;
 wire \fifo0.fifo_store[107][2] ;
 wire \fifo0.fifo_store[107][3] ;
 wire \fifo0.fifo_store[107][4] ;
 wire \fifo0.fifo_store[107][5] ;
 wire \fifo0.fifo_store[107][6] ;
 wire \fifo0.fifo_store[107][7] ;
 wire \fifo0.fifo_store[107][8] ;
 wire \fifo0.fifo_store[107][9] ;
 wire \fifo0.fifo_store[108][0] ;
 wire \fifo0.fifo_store[108][10] ;
 wire \fifo0.fifo_store[108][11] ;
 wire \fifo0.fifo_store[108][12] ;
 wire \fifo0.fifo_store[108][13] ;
 wire \fifo0.fifo_store[108][14] ;
 wire \fifo0.fifo_store[108][15] ;
 wire \fifo0.fifo_store[108][1] ;
 wire \fifo0.fifo_store[108][2] ;
 wire \fifo0.fifo_store[108][3] ;
 wire \fifo0.fifo_store[108][4] ;
 wire \fifo0.fifo_store[108][5] ;
 wire \fifo0.fifo_store[108][6] ;
 wire \fifo0.fifo_store[108][7] ;
 wire \fifo0.fifo_store[108][8] ;
 wire \fifo0.fifo_store[108][9] ;
 wire \fifo0.fifo_store[109][0] ;
 wire \fifo0.fifo_store[109][10] ;
 wire \fifo0.fifo_store[109][11] ;
 wire \fifo0.fifo_store[109][12] ;
 wire \fifo0.fifo_store[109][13] ;
 wire \fifo0.fifo_store[109][14] ;
 wire \fifo0.fifo_store[109][15] ;
 wire \fifo0.fifo_store[109][1] ;
 wire \fifo0.fifo_store[109][2] ;
 wire \fifo0.fifo_store[109][3] ;
 wire \fifo0.fifo_store[109][4] ;
 wire \fifo0.fifo_store[109][5] ;
 wire \fifo0.fifo_store[109][6] ;
 wire \fifo0.fifo_store[109][7] ;
 wire \fifo0.fifo_store[109][8] ;
 wire \fifo0.fifo_store[109][9] ;
 wire \fifo0.fifo_store[10][0] ;
 wire \fifo0.fifo_store[10][10] ;
 wire \fifo0.fifo_store[10][11] ;
 wire \fifo0.fifo_store[10][12] ;
 wire \fifo0.fifo_store[10][13] ;
 wire \fifo0.fifo_store[10][14] ;
 wire \fifo0.fifo_store[10][15] ;
 wire \fifo0.fifo_store[10][1] ;
 wire \fifo0.fifo_store[10][2] ;
 wire \fifo0.fifo_store[10][3] ;
 wire \fifo0.fifo_store[10][4] ;
 wire \fifo0.fifo_store[10][5] ;
 wire \fifo0.fifo_store[10][6] ;
 wire \fifo0.fifo_store[10][7] ;
 wire \fifo0.fifo_store[10][8] ;
 wire \fifo0.fifo_store[10][9] ;
 wire \fifo0.fifo_store[110][0] ;
 wire \fifo0.fifo_store[110][10] ;
 wire \fifo0.fifo_store[110][11] ;
 wire \fifo0.fifo_store[110][12] ;
 wire \fifo0.fifo_store[110][13] ;
 wire \fifo0.fifo_store[110][14] ;
 wire \fifo0.fifo_store[110][15] ;
 wire \fifo0.fifo_store[110][1] ;
 wire \fifo0.fifo_store[110][2] ;
 wire \fifo0.fifo_store[110][3] ;
 wire \fifo0.fifo_store[110][4] ;
 wire \fifo0.fifo_store[110][5] ;
 wire \fifo0.fifo_store[110][6] ;
 wire \fifo0.fifo_store[110][7] ;
 wire \fifo0.fifo_store[110][8] ;
 wire \fifo0.fifo_store[110][9] ;
 wire \fifo0.fifo_store[111][0] ;
 wire \fifo0.fifo_store[111][10] ;
 wire \fifo0.fifo_store[111][11] ;
 wire \fifo0.fifo_store[111][12] ;
 wire \fifo0.fifo_store[111][13] ;
 wire \fifo0.fifo_store[111][14] ;
 wire \fifo0.fifo_store[111][15] ;
 wire \fifo0.fifo_store[111][1] ;
 wire \fifo0.fifo_store[111][2] ;
 wire \fifo0.fifo_store[111][3] ;
 wire \fifo0.fifo_store[111][4] ;
 wire \fifo0.fifo_store[111][5] ;
 wire \fifo0.fifo_store[111][6] ;
 wire \fifo0.fifo_store[111][7] ;
 wire \fifo0.fifo_store[111][8] ;
 wire \fifo0.fifo_store[111][9] ;
 wire \fifo0.fifo_store[112][0] ;
 wire \fifo0.fifo_store[112][10] ;
 wire \fifo0.fifo_store[112][11] ;
 wire \fifo0.fifo_store[112][12] ;
 wire \fifo0.fifo_store[112][13] ;
 wire \fifo0.fifo_store[112][14] ;
 wire \fifo0.fifo_store[112][15] ;
 wire \fifo0.fifo_store[112][1] ;
 wire \fifo0.fifo_store[112][2] ;
 wire \fifo0.fifo_store[112][3] ;
 wire \fifo0.fifo_store[112][4] ;
 wire \fifo0.fifo_store[112][5] ;
 wire \fifo0.fifo_store[112][6] ;
 wire \fifo0.fifo_store[112][7] ;
 wire \fifo0.fifo_store[112][8] ;
 wire \fifo0.fifo_store[112][9] ;
 wire \fifo0.fifo_store[113][0] ;
 wire \fifo0.fifo_store[113][10] ;
 wire \fifo0.fifo_store[113][11] ;
 wire \fifo0.fifo_store[113][12] ;
 wire \fifo0.fifo_store[113][13] ;
 wire \fifo0.fifo_store[113][14] ;
 wire \fifo0.fifo_store[113][15] ;
 wire \fifo0.fifo_store[113][1] ;
 wire \fifo0.fifo_store[113][2] ;
 wire \fifo0.fifo_store[113][3] ;
 wire \fifo0.fifo_store[113][4] ;
 wire \fifo0.fifo_store[113][5] ;
 wire \fifo0.fifo_store[113][6] ;
 wire \fifo0.fifo_store[113][7] ;
 wire \fifo0.fifo_store[113][8] ;
 wire \fifo0.fifo_store[113][9] ;
 wire \fifo0.fifo_store[114][0] ;
 wire \fifo0.fifo_store[114][10] ;
 wire \fifo0.fifo_store[114][11] ;
 wire \fifo0.fifo_store[114][12] ;
 wire \fifo0.fifo_store[114][13] ;
 wire \fifo0.fifo_store[114][14] ;
 wire \fifo0.fifo_store[114][15] ;
 wire \fifo0.fifo_store[114][1] ;
 wire \fifo0.fifo_store[114][2] ;
 wire \fifo0.fifo_store[114][3] ;
 wire \fifo0.fifo_store[114][4] ;
 wire \fifo0.fifo_store[114][5] ;
 wire \fifo0.fifo_store[114][6] ;
 wire \fifo0.fifo_store[114][7] ;
 wire \fifo0.fifo_store[114][8] ;
 wire \fifo0.fifo_store[114][9] ;
 wire \fifo0.fifo_store[115][0] ;
 wire \fifo0.fifo_store[115][10] ;
 wire \fifo0.fifo_store[115][11] ;
 wire \fifo0.fifo_store[115][12] ;
 wire \fifo0.fifo_store[115][13] ;
 wire \fifo0.fifo_store[115][14] ;
 wire \fifo0.fifo_store[115][15] ;
 wire \fifo0.fifo_store[115][1] ;
 wire \fifo0.fifo_store[115][2] ;
 wire \fifo0.fifo_store[115][3] ;
 wire \fifo0.fifo_store[115][4] ;
 wire \fifo0.fifo_store[115][5] ;
 wire \fifo0.fifo_store[115][6] ;
 wire \fifo0.fifo_store[115][7] ;
 wire \fifo0.fifo_store[115][8] ;
 wire \fifo0.fifo_store[115][9] ;
 wire \fifo0.fifo_store[116][0] ;
 wire \fifo0.fifo_store[116][10] ;
 wire \fifo0.fifo_store[116][11] ;
 wire \fifo0.fifo_store[116][12] ;
 wire \fifo0.fifo_store[116][13] ;
 wire \fifo0.fifo_store[116][14] ;
 wire \fifo0.fifo_store[116][15] ;
 wire \fifo0.fifo_store[116][1] ;
 wire \fifo0.fifo_store[116][2] ;
 wire \fifo0.fifo_store[116][3] ;
 wire \fifo0.fifo_store[116][4] ;
 wire \fifo0.fifo_store[116][5] ;
 wire \fifo0.fifo_store[116][6] ;
 wire \fifo0.fifo_store[116][7] ;
 wire \fifo0.fifo_store[116][8] ;
 wire \fifo0.fifo_store[116][9] ;
 wire \fifo0.fifo_store[117][0] ;
 wire \fifo0.fifo_store[117][10] ;
 wire \fifo0.fifo_store[117][11] ;
 wire \fifo0.fifo_store[117][12] ;
 wire \fifo0.fifo_store[117][13] ;
 wire \fifo0.fifo_store[117][14] ;
 wire \fifo0.fifo_store[117][15] ;
 wire \fifo0.fifo_store[117][1] ;
 wire \fifo0.fifo_store[117][2] ;
 wire \fifo0.fifo_store[117][3] ;
 wire \fifo0.fifo_store[117][4] ;
 wire \fifo0.fifo_store[117][5] ;
 wire \fifo0.fifo_store[117][6] ;
 wire \fifo0.fifo_store[117][7] ;
 wire \fifo0.fifo_store[117][8] ;
 wire \fifo0.fifo_store[117][9] ;
 wire \fifo0.fifo_store[118][0] ;
 wire \fifo0.fifo_store[118][10] ;
 wire \fifo0.fifo_store[118][11] ;
 wire \fifo0.fifo_store[118][12] ;
 wire \fifo0.fifo_store[118][13] ;
 wire \fifo0.fifo_store[118][14] ;
 wire \fifo0.fifo_store[118][15] ;
 wire \fifo0.fifo_store[118][1] ;
 wire \fifo0.fifo_store[118][2] ;
 wire \fifo0.fifo_store[118][3] ;
 wire \fifo0.fifo_store[118][4] ;
 wire \fifo0.fifo_store[118][5] ;
 wire \fifo0.fifo_store[118][6] ;
 wire \fifo0.fifo_store[118][7] ;
 wire \fifo0.fifo_store[118][8] ;
 wire \fifo0.fifo_store[118][9] ;
 wire \fifo0.fifo_store[119][0] ;
 wire \fifo0.fifo_store[119][10] ;
 wire \fifo0.fifo_store[119][11] ;
 wire \fifo0.fifo_store[119][12] ;
 wire \fifo0.fifo_store[119][13] ;
 wire \fifo0.fifo_store[119][14] ;
 wire \fifo0.fifo_store[119][15] ;
 wire \fifo0.fifo_store[119][1] ;
 wire \fifo0.fifo_store[119][2] ;
 wire \fifo0.fifo_store[119][3] ;
 wire \fifo0.fifo_store[119][4] ;
 wire \fifo0.fifo_store[119][5] ;
 wire \fifo0.fifo_store[119][6] ;
 wire \fifo0.fifo_store[119][7] ;
 wire \fifo0.fifo_store[119][8] ;
 wire \fifo0.fifo_store[119][9] ;
 wire \fifo0.fifo_store[11][0] ;
 wire \fifo0.fifo_store[11][10] ;
 wire \fifo0.fifo_store[11][11] ;
 wire \fifo0.fifo_store[11][12] ;
 wire \fifo0.fifo_store[11][13] ;
 wire \fifo0.fifo_store[11][14] ;
 wire \fifo0.fifo_store[11][15] ;
 wire \fifo0.fifo_store[11][1] ;
 wire \fifo0.fifo_store[11][2] ;
 wire \fifo0.fifo_store[11][3] ;
 wire \fifo0.fifo_store[11][4] ;
 wire \fifo0.fifo_store[11][5] ;
 wire \fifo0.fifo_store[11][6] ;
 wire \fifo0.fifo_store[11][7] ;
 wire \fifo0.fifo_store[11][8] ;
 wire \fifo0.fifo_store[11][9] ;
 wire \fifo0.fifo_store[120][0] ;
 wire \fifo0.fifo_store[120][10] ;
 wire \fifo0.fifo_store[120][11] ;
 wire \fifo0.fifo_store[120][12] ;
 wire \fifo0.fifo_store[120][13] ;
 wire \fifo0.fifo_store[120][14] ;
 wire \fifo0.fifo_store[120][15] ;
 wire \fifo0.fifo_store[120][1] ;
 wire \fifo0.fifo_store[120][2] ;
 wire \fifo0.fifo_store[120][3] ;
 wire \fifo0.fifo_store[120][4] ;
 wire \fifo0.fifo_store[120][5] ;
 wire \fifo0.fifo_store[120][6] ;
 wire \fifo0.fifo_store[120][7] ;
 wire \fifo0.fifo_store[120][8] ;
 wire \fifo0.fifo_store[120][9] ;
 wire \fifo0.fifo_store[121][0] ;
 wire \fifo0.fifo_store[121][10] ;
 wire \fifo0.fifo_store[121][11] ;
 wire \fifo0.fifo_store[121][12] ;
 wire \fifo0.fifo_store[121][13] ;
 wire \fifo0.fifo_store[121][14] ;
 wire \fifo0.fifo_store[121][15] ;
 wire \fifo0.fifo_store[121][1] ;
 wire \fifo0.fifo_store[121][2] ;
 wire \fifo0.fifo_store[121][3] ;
 wire \fifo0.fifo_store[121][4] ;
 wire \fifo0.fifo_store[121][5] ;
 wire \fifo0.fifo_store[121][6] ;
 wire \fifo0.fifo_store[121][7] ;
 wire \fifo0.fifo_store[121][8] ;
 wire \fifo0.fifo_store[121][9] ;
 wire \fifo0.fifo_store[122][0] ;
 wire \fifo0.fifo_store[122][10] ;
 wire \fifo0.fifo_store[122][11] ;
 wire \fifo0.fifo_store[122][12] ;
 wire \fifo0.fifo_store[122][13] ;
 wire \fifo0.fifo_store[122][14] ;
 wire \fifo0.fifo_store[122][15] ;
 wire \fifo0.fifo_store[122][1] ;
 wire \fifo0.fifo_store[122][2] ;
 wire \fifo0.fifo_store[122][3] ;
 wire \fifo0.fifo_store[122][4] ;
 wire \fifo0.fifo_store[122][5] ;
 wire \fifo0.fifo_store[122][6] ;
 wire \fifo0.fifo_store[122][7] ;
 wire \fifo0.fifo_store[122][8] ;
 wire \fifo0.fifo_store[122][9] ;
 wire \fifo0.fifo_store[123][0] ;
 wire \fifo0.fifo_store[123][10] ;
 wire \fifo0.fifo_store[123][11] ;
 wire \fifo0.fifo_store[123][12] ;
 wire \fifo0.fifo_store[123][13] ;
 wire \fifo0.fifo_store[123][14] ;
 wire \fifo0.fifo_store[123][15] ;
 wire \fifo0.fifo_store[123][1] ;
 wire \fifo0.fifo_store[123][2] ;
 wire \fifo0.fifo_store[123][3] ;
 wire \fifo0.fifo_store[123][4] ;
 wire \fifo0.fifo_store[123][5] ;
 wire \fifo0.fifo_store[123][6] ;
 wire \fifo0.fifo_store[123][7] ;
 wire \fifo0.fifo_store[123][8] ;
 wire \fifo0.fifo_store[123][9] ;
 wire \fifo0.fifo_store[124][0] ;
 wire \fifo0.fifo_store[124][10] ;
 wire \fifo0.fifo_store[124][11] ;
 wire \fifo0.fifo_store[124][12] ;
 wire \fifo0.fifo_store[124][13] ;
 wire \fifo0.fifo_store[124][14] ;
 wire \fifo0.fifo_store[124][15] ;
 wire \fifo0.fifo_store[124][1] ;
 wire \fifo0.fifo_store[124][2] ;
 wire \fifo0.fifo_store[124][3] ;
 wire \fifo0.fifo_store[124][4] ;
 wire \fifo0.fifo_store[124][5] ;
 wire \fifo0.fifo_store[124][6] ;
 wire \fifo0.fifo_store[124][7] ;
 wire \fifo0.fifo_store[124][8] ;
 wire \fifo0.fifo_store[124][9] ;
 wire \fifo0.fifo_store[125][0] ;
 wire \fifo0.fifo_store[125][10] ;
 wire \fifo0.fifo_store[125][11] ;
 wire \fifo0.fifo_store[125][12] ;
 wire \fifo0.fifo_store[125][13] ;
 wire \fifo0.fifo_store[125][14] ;
 wire \fifo0.fifo_store[125][15] ;
 wire \fifo0.fifo_store[125][1] ;
 wire \fifo0.fifo_store[125][2] ;
 wire \fifo0.fifo_store[125][3] ;
 wire \fifo0.fifo_store[125][4] ;
 wire \fifo0.fifo_store[125][5] ;
 wire \fifo0.fifo_store[125][6] ;
 wire \fifo0.fifo_store[125][7] ;
 wire \fifo0.fifo_store[125][8] ;
 wire \fifo0.fifo_store[125][9] ;
 wire \fifo0.fifo_store[126][0] ;
 wire \fifo0.fifo_store[126][10] ;
 wire \fifo0.fifo_store[126][11] ;
 wire \fifo0.fifo_store[126][12] ;
 wire \fifo0.fifo_store[126][13] ;
 wire \fifo0.fifo_store[126][14] ;
 wire \fifo0.fifo_store[126][15] ;
 wire \fifo0.fifo_store[126][1] ;
 wire \fifo0.fifo_store[126][2] ;
 wire \fifo0.fifo_store[126][3] ;
 wire \fifo0.fifo_store[126][4] ;
 wire \fifo0.fifo_store[126][5] ;
 wire \fifo0.fifo_store[126][6] ;
 wire \fifo0.fifo_store[126][7] ;
 wire \fifo0.fifo_store[126][8] ;
 wire \fifo0.fifo_store[126][9] ;
 wire \fifo0.fifo_store[127][0] ;
 wire \fifo0.fifo_store[127][10] ;
 wire \fifo0.fifo_store[127][11] ;
 wire \fifo0.fifo_store[127][12] ;
 wire \fifo0.fifo_store[127][13] ;
 wire \fifo0.fifo_store[127][14] ;
 wire \fifo0.fifo_store[127][15] ;
 wire \fifo0.fifo_store[127][1] ;
 wire \fifo0.fifo_store[127][2] ;
 wire \fifo0.fifo_store[127][3] ;
 wire \fifo0.fifo_store[127][4] ;
 wire \fifo0.fifo_store[127][5] ;
 wire \fifo0.fifo_store[127][6] ;
 wire \fifo0.fifo_store[127][7] ;
 wire \fifo0.fifo_store[127][8] ;
 wire \fifo0.fifo_store[127][9] ;
 wire \fifo0.fifo_store[12][0] ;
 wire \fifo0.fifo_store[12][10] ;
 wire \fifo0.fifo_store[12][11] ;
 wire \fifo0.fifo_store[12][12] ;
 wire \fifo0.fifo_store[12][13] ;
 wire \fifo0.fifo_store[12][14] ;
 wire \fifo0.fifo_store[12][15] ;
 wire \fifo0.fifo_store[12][1] ;
 wire \fifo0.fifo_store[12][2] ;
 wire \fifo0.fifo_store[12][3] ;
 wire \fifo0.fifo_store[12][4] ;
 wire \fifo0.fifo_store[12][5] ;
 wire \fifo0.fifo_store[12][6] ;
 wire \fifo0.fifo_store[12][7] ;
 wire \fifo0.fifo_store[12][8] ;
 wire \fifo0.fifo_store[12][9] ;
 wire \fifo0.fifo_store[13][0] ;
 wire \fifo0.fifo_store[13][10] ;
 wire \fifo0.fifo_store[13][11] ;
 wire \fifo0.fifo_store[13][12] ;
 wire \fifo0.fifo_store[13][13] ;
 wire \fifo0.fifo_store[13][14] ;
 wire \fifo0.fifo_store[13][15] ;
 wire \fifo0.fifo_store[13][1] ;
 wire \fifo0.fifo_store[13][2] ;
 wire \fifo0.fifo_store[13][3] ;
 wire \fifo0.fifo_store[13][4] ;
 wire \fifo0.fifo_store[13][5] ;
 wire \fifo0.fifo_store[13][6] ;
 wire \fifo0.fifo_store[13][7] ;
 wire \fifo0.fifo_store[13][8] ;
 wire \fifo0.fifo_store[13][9] ;
 wire \fifo0.fifo_store[14][0] ;
 wire \fifo0.fifo_store[14][10] ;
 wire \fifo0.fifo_store[14][11] ;
 wire \fifo0.fifo_store[14][12] ;
 wire \fifo0.fifo_store[14][13] ;
 wire \fifo0.fifo_store[14][14] ;
 wire \fifo0.fifo_store[14][15] ;
 wire \fifo0.fifo_store[14][1] ;
 wire \fifo0.fifo_store[14][2] ;
 wire \fifo0.fifo_store[14][3] ;
 wire \fifo0.fifo_store[14][4] ;
 wire \fifo0.fifo_store[14][5] ;
 wire \fifo0.fifo_store[14][6] ;
 wire \fifo0.fifo_store[14][7] ;
 wire \fifo0.fifo_store[14][8] ;
 wire \fifo0.fifo_store[14][9] ;
 wire \fifo0.fifo_store[15][0] ;
 wire \fifo0.fifo_store[15][10] ;
 wire \fifo0.fifo_store[15][11] ;
 wire \fifo0.fifo_store[15][12] ;
 wire \fifo0.fifo_store[15][13] ;
 wire \fifo0.fifo_store[15][14] ;
 wire \fifo0.fifo_store[15][15] ;
 wire \fifo0.fifo_store[15][1] ;
 wire \fifo0.fifo_store[15][2] ;
 wire \fifo0.fifo_store[15][3] ;
 wire \fifo0.fifo_store[15][4] ;
 wire \fifo0.fifo_store[15][5] ;
 wire \fifo0.fifo_store[15][6] ;
 wire \fifo0.fifo_store[15][7] ;
 wire \fifo0.fifo_store[15][8] ;
 wire \fifo0.fifo_store[15][9] ;
 wire \fifo0.fifo_store[16][0] ;
 wire \fifo0.fifo_store[16][10] ;
 wire \fifo0.fifo_store[16][11] ;
 wire \fifo0.fifo_store[16][12] ;
 wire \fifo0.fifo_store[16][13] ;
 wire \fifo0.fifo_store[16][14] ;
 wire \fifo0.fifo_store[16][15] ;
 wire \fifo0.fifo_store[16][1] ;
 wire \fifo0.fifo_store[16][2] ;
 wire \fifo0.fifo_store[16][3] ;
 wire \fifo0.fifo_store[16][4] ;
 wire \fifo0.fifo_store[16][5] ;
 wire \fifo0.fifo_store[16][6] ;
 wire \fifo0.fifo_store[16][7] ;
 wire \fifo0.fifo_store[16][8] ;
 wire \fifo0.fifo_store[16][9] ;
 wire \fifo0.fifo_store[17][0] ;
 wire \fifo0.fifo_store[17][10] ;
 wire \fifo0.fifo_store[17][11] ;
 wire \fifo0.fifo_store[17][12] ;
 wire \fifo0.fifo_store[17][13] ;
 wire \fifo0.fifo_store[17][14] ;
 wire \fifo0.fifo_store[17][15] ;
 wire \fifo0.fifo_store[17][1] ;
 wire \fifo0.fifo_store[17][2] ;
 wire \fifo0.fifo_store[17][3] ;
 wire \fifo0.fifo_store[17][4] ;
 wire \fifo0.fifo_store[17][5] ;
 wire \fifo0.fifo_store[17][6] ;
 wire \fifo0.fifo_store[17][7] ;
 wire \fifo0.fifo_store[17][8] ;
 wire \fifo0.fifo_store[17][9] ;
 wire \fifo0.fifo_store[18][0] ;
 wire \fifo0.fifo_store[18][10] ;
 wire \fifo0.fifo_store[18][11] ;
 wire \fifo0.fifo_store[18][12] ;
 wire \fifo0.fifo_store[18][13] ;
 wire \fifo0.fifo_store[18][14] ;
 wire \fifo0.fifo_store[18][15] ;
 wire \fifo0.fifo_store[18][1] ;
 wire \fifo0.fifo_store[18][2] ;
 wire \fifo0.fifo_store[18][3] ;
 wire \fifo0.fifo_store[18][4] ;
 wire \fifo0.fifo_store[18][5] ;
 wire \fifo0.fifo_store[18][6] ;
 wire \fifo0.fifo_store[18][7] ;
 wire \fifo0.fifo_store[18][8] ;
 wire \fifo0.fifo_store[18][9] ;
 wire \fifo0.fifo_store[19][0] ;
 wire \fifo0.fifo_store[19][10] ;
 wire \fifo0.fifo_store[19][11] ;
 wire \fifo0.fifo_store[19][12] ;
 wire \fifo0.fifo_store[19][13] ;
 wire \fifo0.fifo_store[19][14] ;
 wire \fifo0.fifo_store[19][15] ;
 wire \fifo0.fifo_store[19][1] ;
 wire \fifo0.fifo_store[19][2] ;
 wire \fifo0.fifo_store[19][3] ;
 wire \fifo0.fifo_store[19][4] ;
 wire \fifo0.fifo_store[19][5] ;
 wire \fifo0.fifo_store[19][6] ;
 wire \fifo0.fifo_store[19][7] ;
 wire \fifo0.fifo_store[19][8] ;
 wire \fifo0.fifo_store[19][9] ;
 wire \fifo0.fifo_store[1][0] ;
 wire \fifo0.fifo_store[1][10] ;
 wire \fifo0.fifo_store[1][11] ;
 wire \fifo0.fifo_store[1][12] ;
 wire \fifo0.fifo_store[1][13] ;
 wire \fifo0.fifo_store[1][14] ;
 wire \fifo0.fifo_store[1][15] ;
 wire \fifo0.fifo_store[1][1] ;
 wire \fifo0.fifo_store[1][2] ;
 wire \fifo0.fifo_store[1][3] ;
 wire \fifo0.fifo_store[1][4] ;
 wire \fifo0.fifo_store[1][5] ;
 wire \fifo0.fifo_store[1][6] ;
 wire \fifo0.fifo_store[1][7] ;
 wire \fifo0.fifo_store[1][8] ;
 wire \fifo0.fifo_store[1][9] ;
 wire \fifo0.fifo_store[20][0] ;
 wire \fifo0.fifo_store[20][10] ;
 wire \fifo0.fifo_store[20][11] ;
 wire \fifo0.fifo_store[20][12] ;
 wire \fifo0.fifo_store[20][13] ;
 wire \fifo0.fifo_store[20][14] ;
 wire \fifo0.fifo_store[20][15] ;
 wire \fifo0.fifo_store[20][1] ;
 wire \fifo0.fifo_store[20][2] ;
 wire \fifo0.fifo_store[20][3] ;
 wire \fifo0.fifo_store[20][4] ;
 wire \fifo0.fifo_store[20][5] ;
 wire \fifo0.fifo_store[20][6] ;
 wire \fifo0.fifo_store[20][7] ;
 wire \fifo0.fifo_store[20][8] ;
 wire \fifo0.fifo_store[20][9] ;
 wire \fifo0.fifo_store[21][0] ;
 wire \fifo0.fifo_store[21][10] ;
 wire \fifo0.fifo_store[21][11] ;
 wire \fifo0.fifo_store[21][12] ;
 wire \fifo0.fifo_store[21][13] ;
 wire \fifo0.fifo_store[21][14] ;
 wire \fifo0.fifo_store[21][15] ;
 wire \fifo0.fifo_store[21][1] ;
 wire \fifo0.fifo_store[21][2] ;
 wire \fifo0.fifo_store[21][3] ;
 wire \fifo0.fifo_store[21][4] ;
 wire \fifo0.fifo_store[21][5] ;
 wire \fifo0.fifo_store[21][6] ;
 wire \fifo0.fifo_store[21][7] ;
 wire \fifo0.fifo_store[21][8] ;
 wire \fifo0.fifo_store[21][9] ;
 wire \fifo0.fifo_store[22][0] ;
 wire \fifo0.fifo_store[22][10] ;
 wire \fifo0.fifo_store[22][11] ;
 wire \fifo0.fifo_store[22][12] ;
 wire \fifo0.fifo_store[22][13] ;
 wire \fifo0.fifo_store[22][14] ;
 wire \fifo0.fifo_store[22][15] ;
 wire \fifo0.fifo_store[22][1] ;
 wire \fifo0.fifo_store[22][2] ;
 wire \fifo0.fifo_store[22][3] ;
 wire \fifo0.fifo_store[22][4] ;
 wire \fifo0.fifo_store[22][5] ;
 wire \fifo0.fifo_store[22][6] ;
 wire \fifo0.fifo_store[22][7] ;
 wire \fifo0.fifo_store[22][8] ;
 wire \fifo0.fifo_store[22][9] ;
 wire \fifo0.fifo_store[23][0] ;
 wire \fifo0.fifo_store[23][10] ;
 wire \fifo0.fifo_store[23][11] ;
 wire \fifo0.fifo_store[23][12] ;
 wire \fifo0.fifo_store[23][13] ;
 wire \fifo0.fifo_store[23][14] ;
 wire \fifo0.fifo_store[23][15] ;
 wire \fifo0.fifo_store[23][1] ;
 wire \fifo0.fifo_store[23][2] ;
 wire \fifo0.fifo_store[23][3] ;
 wire \fifo0.fifo_store[23][4] ;
 wire \fifo0.fifo_store[23][5] ;
 wire \fifo0.fifo_store[23][6] ;
 wire \fifo0.fifo_store[23][7] ;
 wire \fifo0.fifo_store[23][8] ;
 wire \fifo0.fifo_store[23][9] ;
 wire \fifo0.fifo_store[24][0] ;
 wire \fifo0.fifo_store[24][10] ;
 wire \fifo0.fifo_store[24][11] ;
 wire \fifo0.fifo_store[24][12] ;
 wire \fifo0.fifo_store[24][13] ;
 wire \fifo0.fifo_store[24][14] ;
 wire \fifo0.fifo_store[24][15] ;
 wire \fifo0.fifo_store[24][1] ;
 wire \fifo0.fifo_store[24][2] ;
 wire \fifo0.fifo_store[24][3] ;
 wire \fifo0.fifo_store[24][4] ;
 wire \fifo0.fifo_store[24][5] ;
 wire \fifo0.fifo_store[24][6] ;
 wire \fifo0.fifo_store[24][7] ;
 wire \fifo0.fifo_store[24][8] ;
 wire \fifo0.fifo_store[24][9] ;
 wire \fifo0.fifo_store[25][0] ;
 wire \fifo0.fifo_store[25][10] ;
 wire \fifo0.fifo_store[25][11] ;
 wire \fifo0.fifo_store[25][12] ;
 wire \fifo0.fifo_store[25][13] ;
 wire \fifo0.fifo_store[25][14] ;
 wire \fifo0.fifo_store[25][15] ;
 wire \fifo0.fifo_store[25][1] ;
 wire \fifo0.fifo_store[25][2] ;
 wire \fifo0.fifo_store[25][3] ;
 wire \fifo0.fifo_store[25][4] ;
 wire \fifo0.fifo_store[25][5] ;
 wire \fifo0.fifo_store[25][6] ;
 wire \fifo0.fifo_store[25][7] ;
 wire \fifo0.fifo_store[25][8] ;
 wire \fifo0.fifo_store[25][9] ;
 wire \fifo0.fifo_store[26][0] ;
 wire \fifo0.fifo_store[26][10] ;
 wire \fifo0.fifo_store[26][11] ;
 wire \fifo0.fifo_store[26][12] ;
 wire \fifo0.fifo_store[26][13] ;
 wire \fifo0.fifo_store[26][14] ;
 wire \fifo0.fifo_store[26][15] ;
 wire \fifo0.fifo_store[26][1] ;
 wire \fifo0.fifo_store[26][2] ;
 wire \fifo0.fifo_store[26][3] ;
 wire \fifo0.fifo_store[26][4] ;
 wire \fifo0.fifo_store[26][5] ;
 wire \fifo0.fifo_store[26][6] ;
 wire \fifo0.fifo_store[26][7] ;
 wire \fifo0.fifo_store[26][8] ;
 wire \fifo0.fifo_store[26][9] ;
 wire \fifo0.fifo_store[27][0] ;
 wire \fifo0.fifo_store[27][10] ;
 wire \fifo0.fifo_store[27][11] ;
 wire \fifo0.fifo_store[27][12] ;
 wire \fifo0.fifo_store[27][13] ;
 wire \fifo0.fifo_store[27][14] ;
 wire \fifo0.fifo_store[27][15] ;
 wire \fifo0.fifo_store[27][1] ;
 wire \fifo0.fifo_store[27][2] ;
 wire \fifo0.fifo_store[27][3] ;
 wire \fifo0.fifo_store[27][4] ;
 wire \fifo0.fifo_store[27][5] ;
 wire \fifo0.fifo_store[27][6] ;
 wire \fifo0.fifo_store[27][7] ;
 wire \fifo0.fifo_store[27][8] ;
 wire \fifo0.fifo_store[27][9] ;
 wire \fifo0.fifo_store[28][0] ;
 wire \fifo0.fifo_store[28][10] ;
 wire \fifo0.fifo_store[28][11] ;
 wire \fifo0.fifo_store[28][12] ;
 wire \fifo0.fifo_store[28][13] ;
 wire \fifo0.fifo_store[28][14] ;
 wire \fifo0.fifo_store[28][15] ;
 wire \fifo0.fifo_store[28][1] ;
 wire \fifo0.fifo_store[28][2] ;
 wire \fifo0.fifo_store[28][3] ;
 wire \fifo0.fifo_store[28][4] ;
 wire \fifo0.fifo_store[28][5] ;
 wire \fifo0.fifo_store[28][6] ;
 wire \fifo0.fifo_store[28][7] ;
 wire \fifo0.fifo_store[28][8] ;
 wire \fifo0.fifo_store[28][9] ;
 wire \fifo0.fifo_store[29][0] ;
 wire \fifo0.fifo_store[29][10] ;
 wire \fifo0.fifo_store[29][11] ;
 wire \fifo0.fifo_store[29][12] ;
 wire \fifo0.fifo_store[29][13] ;
 wire \fifo0.fifo_store[29][14] ;
 wire \fifo0.fifo_store[29][15] ;
 wire \fifo0.fifo_store[29][1] ;
 wire \fifo0.fifo_store[29][2] ;
 wire \fifo0.fifo_store[29][3] ;
 wire \fifo0.fifo_store[29][4] ;
 wire \fifo0.fifo_store[29][5] ;
 wire \fifo0.fifo_store[29][6] ;
 wire \fifo0.fifo_store[29][7] ;
 wire \fifo0.fifo_store[29][8] ;
 wire \fifo0.fifo_store[29][9] ;
 wire \fifo0.fifo_store[2][0] ;
 wire \fifo0.fifo_store[2][10] ;
 wire \fifo0.fifo_store[2][11] ;
 wire \fifo0.fifo_store[2][12] ;
 wire \fifo0.fifo_store[2][13] ;
 wire \fifo0.fifo_store[2][14] ;
 wire \fifo0.fifo_store[2][15] ;
 wire \fifo0.fifo_store[2][1] ;
 wire \fifo0.fifo_store[2][2] ;
 wire \fifo0.fifo_store[2][3] ;
 wire \fifo0.fifo_store[2][4] ;
 wire \fifo0.fifo_store[2][5] ;
 wire \fifo0.fifo_store[2][6] ;
 wire \fifo0.fifo_store[2][7] ;
 wire \fifo0.fifo_store[2][8] ;
 wire \fifo0.fifo_store[2][9] ;
 wire \fifo0.fifo_store[30][0] ;
 wire \fifo0.fifo_store[30][10] ;
 wire \fifo0.fifo_store[30][11] ;
 wire \fifo0.fifo_store[30][12] ;
 wire \fifo0.fifo_store[30][13] ;
 wire \fifo0.fifo_store[30][14] ;
 wire \fifo0.fifo_store[30][15] ;
 wire \fifo0.fifo_store[30][1] ;
 wire \fifo0.fifo_store[30][2] ;
 wire \fifo0.fifo_store[30][3] ;
 wire \fifo0.fifo_store[30][4] ;
 wire \fifo0.fifo_store[30][5] ;
 wire \fifo0.fifo_store[30][6] ;
 wire \fifo0.fifo_store[30][7] ;
 wire \fifo0.fifo_store[30][8] ;
 wire \fifo0.fifo_store[30][9] ;
 wire \fifo0.fifo_store[31][0] ;
 wire \fifo0.fifo_store[31][10] ;
 wire \fifo0.fifo_store[31][11] ;
 wire \fifo0.fifo_store[31][12] ;
 wire \fifo0.fifo_store[31][13] ;
 wire \fifo0.fifo_store[31][14] ;
 wire \fifo0.fifo_store[31][15] ;
 wire \fifo0.fifo_store[31][1] ;
 wire \fifo0.fifo_store[31][2] ;
 wire \fifo0.fifo_store[31][3] ;
 wire \fifo0.fifo_store[31][4] ;
 wire \fifo0.fifo_store[31][5] ;
 wire \fifo0.fifo_store[31][6] ;
 wire \fifo0.fifo_store[31][7] ;
 wire \fifo0.fifo_store[31][8] ;
 wire \fifo0.fifo_store[31][9] ;
 wire \fifo0.fifo_store[32][0] ;
 wire \fifo0.fifo_store[32][10] ;
 wire \fifo0.fifo_store[32][11] ;
 wire \fifo0.fifo_store[32][12] ;
 wire \fifo0.fifo_store[32][13] ;
 wire \fifo0.fifo_store[32][14] ;
 wire \fifo0.fifo_store[32][15] ;
 wire \fifo0.fifo_store[32][1] ;
 wire \fifo0.fifo_store[32][2] ;
 wire \fifo0.fifo_store[32][3] ;
 wire \fifo0.fifo_store[32][4] ;
 wire \fifo0.fifo_store[32][5] ;
 wire \fifo0.fifo_store[32][6] ;
 wire \fifo0.fifo_store[32][7] ;
 wire \fifo0.fifo_store[32][8] ;
 wire \fifo0.fifo_store[32][9] ;
 wire \fifo0.fifo_store[33][0] ;
 wire \fifo0.fifo_store[33][10] ;
 wire \fifo0.fifo_store[33][11] ;
 wire \fifo0.fifo_store[33][12] ;
 wire \fifo0.fifo_store[33][13] ;
 wire \fifo0.fifo_store[33][14] ;
 wire \fifo0.fifo_store[33][15] ;
 wire \fifo0.fifo_store[33][1] ;
 wire \fifo0.fifo_store[33][2] ;
 wire \fifo0.fifo_store[33][3] ;
 wire \fifo0.fifo_store[33][4] ;
 wire \fifo0.fifo_store[33][5] ;
 wire \fifo0.fifo_store[33][6] ;
 wire \fifo0.fifo_store[33][7] ;
 wire \fifo0.fifo_store[33][8] ;
 wire \fifo0.fifo_store[33][9] ;
 wire \fifo0.fifo_store[34][0] ;
 wire \fifo0.fifo_store[34][10] ;
 wire \fifo0.fifo_store[34][11] ;
 wire \fifo0.fifo_store[34][12] ;
 wire \fifo0.fifo_store[34][13] ;
 wire \fifo0.fifo_store[34][14] ;
 wire \fifo0.fifo_store[34][15] ;
 wire \fifo0.fifo_store[34][1] ;
 wire \fifo0.fifo_store[34][2] ;
 wire \fifo0.fifo_store[34][3] ;
 wire \fifo0.fifo_store[34][4] ;
 wire \fifo0.fifo_store[34][5] ;
 wire \fifo0.fifo_store[34][6] ;
 wire \fifo0.fifo_store[34][7] ;
 wire \fifo0.fifo_store[34][8] ;
 wire \fifo0.fifo_store[34][9] ;
 wire \fifo0.fifo_store[35][0] ;
 wire \fifo0.fifo_store[35][10] ;
 wire \fifo0.fifo_store[35][11] ;
 wire \fifo0.fifo_store[35][12] ;
 wire \fifo0.fifo_store[35][13] ;
 wire \fifo0.fifo_store[35][14] ;
 wire \fifo0.fifo_store[35][15] ;
 wire \fifo0.fifo_store[35][1] ;
 wire \fifo0.fifo_store[35][2] ;
 wire \fifo0.fifo_store[35][3] ;
 wire \fifo0.fifo_store[35][4] ;
 wire \fifo0.fifo_store[35][5] ;
 wire \fifo0.fifo_store[35][6] ;
 wire \fifo0.fifo_store[35][7] ;
 wire \fifo0.fifo_store[35][8] ;
 wire \fifo0.fifo_store[35][9] ;
 wire \fifo0.fifo_store[36][0] ;
 wire \fifo0.fifo_store[36][10] ;
 wire \fifo0.fifo_store[36][11] ;
 wire \fifo0.fifo_store[36][12] ;
 wire \fifo0.fifo_store[36][13] ;
 wire \fifo0.fifo_store[36][14] ;
 wire \fifo0.fifo_store[36][15] ;
 wire \fifo0.fifo_store[36][1] ;
 wire \fifo0.fifo_store[36][2] ;
 wire \fifo0.fifo_store[36][3] ;
 wire \fifo0.fifo_store[36][4] ;
 wire \fifo0.fifo_store[36][5] ;
 wire \fifo0.fifo_store[36][6] ;
 wire \fifo0.fifo_store[36][7] ;
 wire \fifo0.fifo_store[36][8] ;
 wire \fifo0.fifo_store[36][9] ;
 wire \fifo0.fifo_store[37][0] ;
 wire \fifo0.fifo_store[37][10] ;
 wire \fifo0.fifo_store[37][11] ;
 wire \fifo0.fifo_store[37][12] ;
 wire \fifo0.fifo_store[37][13] ;
 wire \fifo0.fifo_store[37][14] ;
 wire \fifo0.fifo_store[37][15] ;
 wire \fifo0.fifo_store[37][1] ;
 wire \fifo0.fifo_store[37][2] ;
 wire \fifo0.fifo_store[37][3] ;
 wire \fifo0.fifo_store[37][4] ;
 wire \fifo0.fifo_store[37][5] ;
 wire \fifo0.fifo_store[37][6] ;
 wire \fifo0.fifo_store[37][7] ;
 wire \fifo0.fifo_store[37][8] ;
 wire \fifo0.fifo_store[37][9] ;
 wire \fifo0.fifo_store[38][0] ;
 wire \fifo0.fifo_store[38][10] ;
 wire \fifo0.fifo_store[38][11] ;
 wire \fifo0.fifo_store[38][12] ;
 wire \fifo0.fifo_store[38][13] ;
 wire \fifo0.fifo_store[38][14] ;
 wire \fifo0.fifo_store[38][15] ;
 wire \fifo0.fifo_store[38][1] ;
 wire \fifo0.fifo_store[38][2] ;
 wire \fifo0.fifo_store[38][3] ;
 wire \fifo0.fifo_store[38][4] ;
 wire \fifo0.fifo_store[38][5] ;
 wire \fifo0.fifo_store[38][6] ;
 wire \fifo0.fifo_store[38][7] ;
 wire \fifo0.fifo_store[38][8] ;
 wire \fifo0.fifo_store[38][9] ;
 wire \fifo0.fifo_store[39][0] ;
 wire \fifo0.fifo_store[39][10] ;
 wire \fifo0.fifo_store[39][11] ;
 wire \fifo0.fifo_store[39][12] ;
 wire \fifo0.fifo_store[39][13] ;
 wire \fifo0.fifo_store[39][14] ;
 wire \fifo0.fifo_store[39][15] ;
 wire \fifo0.fifo_store[39][1] ;
 wire \fifo0.fifo_store[39][2] ;
 wire \fifo0.fifo_store[39][3] ;
 wire \fifo0.fifo_store[39][4] ;
 wire \fifo0.fifo_store[39][5] ;
 wire \fifo0.fifo_store[39][6] ;
 wire \fifo0.fifo_store[39][7] ;
 wire \fifo0.fifo_store[39][8] ;
 wire \fifo0.fifo_store[39][9] ;
 wire \fifo0.fifo_store[3][0] ;
 wire \fifo0.fifo_store[3][10] ;
 wire \fifo0.fifo_store[3][11] ;
 wire \fifo0.fifo_store[3][12] ;
 wire \fifo0.fifo_store[3][13] ;
 wire \fifo0.fifo_store[3][14] ;
 wire \fifo0.fifo_store[3][15] ;
 wire \fifo0.fifo_store[3][1] ;
 wire \fifo0.fifo_store[3][2] ;
 wire \fifo0.fifo_store[3][3] ;
 wire \fifo0.fifo_store[3][4] ;
 wire \fifo0.fifo_store[3][5] ;
 wire \fifo0.fifo_store[3][6] ;
 wire \fifo0.fifo_store[3][7] ;
 wire \fifo0.fifo_store[3][8] ;
 wire \fifo0.fifo_store[3][9] ;
 wire \fifo0.fifo_store[40][0] ;
 wire \fifo0.fifo_store[40][10] ;
 wire \fifo0.fifo_store[40][11] ;
 wire \fifo0.fifo_store[40][12] ;
 wire \fifo0.fifo_store[40][13] ;
 wire \fifo0.fifo_store[40][14] ;
 wire \fifo0.fifo_store[40][15] ;
 wire \fifo0.fifo_store[40][1] ;
 wire \fifo0.fifo_store[40][2] ;
 wire \fifo0.fifo_store[40][3] ;
 wire \fifo0.fifo_store[40][4] ;
 wire \fifo0.fifo_store[40][5] ;
 wire \fifo0.fifo_store[40][6] ;
 wire \fifo0.fifo_store[40][7] ;
 wire \fifo0.fifo_store[40][8] ;
 wire \fifo0.fifo_store[40][9] ;
 wire \fifo0.fifo_store[41][0] ;
 wire \fifo0.fifo_store[41][10] ;
 wire \fifo0.fifo_store[41][11] ;
 wire \fifo0.fifo_store[41][12] ;
 wire \fifo0.fifo_store[41][13] ;
 wire \fifo0.fifo_store[41][14] ;
 wire \fifo0.fifo_store[41][15] ;
 wire \fifo0.fifo_store[41][1] ;
 wire \fifo0.fifo_store[41][2] ;
 wire \fifo0.fifo_store[41][3] ;
 wire \fifo0.fifo_store[41][4] ;
 wire \fifo0.fifo_store[41][5] ;
 wire \fifo0.fifo_store[41][6] ;
 wire \fifo0.fifo_store[41][7] ;
 wire \fifo0.fifo_store[41][8] ;
 wire \fifo0.fifo_store[41][9] ;
 wire \fifo0.fifo_store[42][0] ;
 wire \fifo0.fifo_store[42][10] ;
 wire \fifo0.fifo_store[42][11] ;
 wire \fifo0.fifo_store[42][12] ;
 wire \fifo0.fifo_store[42][13] ;
 wire \fifo0.fifo_store[42][14] ;
 wire \fifo0.fifo_store[42][15] ;
 wire \fifo0.fifo_store[42][1] ;
 wire \fifo0.fifo_store[42][2] ;
 wire \fifo0.fifo_store[42][3] ;
 wire \fifo0.fifo_store[42][4] ;
 wire \fifo0.fifo_store[42][5] ;
 wire \fifo0.fifo_store[42][6] ;
 wire \fifo0.fifo_store[42][7] ;
 wire \fifo0.fifo_store[42][8] ;
 wire \fifo0.fifo_store[42][9] ;
 wire \fifo0.fifo_store[43][0] ;
 wire \fifo0.fifo_store[43][10] ;
 wire \fifo0.fifo_store[43][11] ;
 wire \fifo0.fifo_store[43][12] ;
 wire \fifo0.fifo_store[43][13] ;
 wire \fifo0.fifo_store[43][14] ;
 wire \fifo0.fifo_store[43][15] ;
 wire \fifo0.fifo_store[43][1] ;
 wire \fifo0.fifo_store[43][2] ;
 wire \fifo0.fifo_store[43][3] ;
 wire \fifo0.fifo_store[43][4] ;
 wire \fifo0.fifo_store[43][5] ;
 wire \fifo0.fifo_store[43][6] ;
 wire \fifo0.fifo_store[43][7] ;
 wire \fifo0.fifo_store[43][8] ;
 wire \fifo0.fifo_store[43][9] ;
 wire \fifo0.fifo_store[44][0] ;
 wire \fifo0.fifo_store[44][10] ;
 wire \fifo0.fifo_store[44][11] ;
 wire \fifo0.fifo_store[44][12] ;
 wire \fifo0.fifo_store[44][13] ;
 wire \fifo0.fifo_store[44][14] ;
 wire \fifo0.fifo_store[44][15] ;
 wire \fifo0.fifo_store[44][1] ;
 wire \fifo0.fifo_store[44][2] ;
 wire \fifo0.fifo_store[44][3] ;
 wire \fifo0.fifo_store[44][4] ;
 wire \fifo0.fifo_store[44][5] ;
 wire \fifo0.fifo_store[44][6] ;
 wire \fifo0.fifo_store[44][7] ;
 wire \fifo0.fifo_store[44][8] ;
 wire \fifo0.fifo_store[44][9] ;
 wire \fifo0.fifo_store[45][0] ;
 wire \fifo0.fifo_store[45][10] ;
 wire \fifo0.fifo_store[45][11] ;
 wire \fifo0.fifo_store[45][12] ;
 wire \fifo0.fifo_store[45][13] ;
 wire \fifo0.fifo_store[45][14] ;
 wire \fifo0.fifo_store[45][15] ;
 wire \fifo0.fifo_store[45][1] ;
 wire \fifo0.fifo_store[45][2] ;
 wire \fifo0.fifo_store[45][3] ;
 wire \fifo0.fifo_store[45][4] ;
 wire \fifo0.fifo_store[45][5] ;
 wire \fifo0.fifo_store[45][6] ;
 wire \fifo0.fifo_store[45][7] ;
 wire \fifo0.fifo_store[45][8] ;
 wire \fifo0.fifo_store[45][9] ;
 wire \fifo0.fifo_store[46][0] ;
 wire \fifo0.fifo_store[46][10] ;
 wire \fifo0.fifo_store[46][11] ;
 wire \fifo0.fifo_store[46][12] ;
 wire \fifo0.fifo_store[46][13] ;
 wire \fifo0.fifo_store[46][14] ;
 wire \fifo0.fifo_store[46][15] ;
 wire \fifo0.fifo_store[46][1] ;
 wire \fifo0.fifo_store[46][2] ;
 wire \fifo0.fifo_store[46][3] ;
 wire \fifo0.fifo_store[46][4] ;
 wire \fifo0.fifo_store[46][5] ;
 wire \fifo0.fifo_store[46][6] ;
 wire \fifo0.fifo_store[46][7] ;
 wire \fifo0.fifo_store[46][8] ;
 wire \fifo0.fifo_store[46][9] ;
 wire \fifo0.fifo_store[47][0] ;
 wire \fifo0.fifo_store[47][10] ;
 wire \fifo0.fifo_store[47][11] ;
 wire \fifo0.fifo_store[47][12] ;
 wire \fifo0.fifo_store[47][13] ;
 wire \fifo0.fifo_store[47][14] ;
 wire \fifo0.fifo_store[47][15] ;
 wire \fifo0.fifo_store[47][1] ;
 wire \fifo0.fifo_store[47][2] ;
 wire \fifo0.fifo_store[47][3] ;
 wire \fifo0.fifo_store[47][4] ;
 wire \fifo0.fifo_store[47][5] ;
 wire \fifo0.fifo_store[47][6] ;
 wire \fifo0.fifo_store[47][7] ;
 wire \fifo0.fifo_store[47][8] ;
 wire \fifo0.fifo_store[47][9] ;
 wire \fifo0.fifo_store[48][0] ;
 wire \fifo0.fifo_store[48][10] ;
 wire \fifo0.fifo_store[48][11] ;
 wire \fifo0.fifo_store[48][12] ;
 wire \fifo0.fifo_store[48][13] ;
 wire \fifo0.fifo_store[48][14] ;
 wire \fifo0.fifo_store[48][15] ;
 wire \fifo0.fifo_store[48][1] ;
 wire \fifo0.fifo_store[48][2] ;
 wire \fifo0.fifo_store[48][3] ;
 wire \fifo0.fifo_store[48][4] ;
 wire \fifo0.fifo_store[48][5] ;
 wire \fifo0.fifo_store[48][6] ;
 wire \fifo0.fifo_store[48][7] ;
 wire \fifo0.fifo_store[48][8] ;
 wire \fifo0.fifo_store[48][9] ;
 wire \fifo0.fifo_store[49][0] ;
 wire \fifo0.fifo_store[49][10] ;
 wire \fifo0.fifo_store[49][11] ;
 wire \fifo0.fifo_store[49][12] ;
 wire \fifo0.fifo_store[49][13] ;
 wire \fifo0.fifo_store[49][14] ;
 wire \fifo0.fifo_store[49][15] ;
 wire \fifo0.fifo_store[49][1] ;
 wire \fifo0.fifo_store[49][2] ;
 wire \fifo0.fifo_store[49][3] ;
 wire \fifo0.fifo_store[49][4] ;
 wire \fifo0.fifo_store[49][5] ;
 wire \fifo0.fifo_store[49][6] ;
 wire \fifo0.fifo_store[49][7] ;
 wire \fifo0.fifo_store[49][8] ;
 wire \fifo0.fifo_store[49][9] ;
 wire \fifo0.fifo_store[4][0] ;
 wire \fifo0.fifo_store[4][10] ;
 wire \fifo0.fifo_store[4][11] ;
 wire \fifo0.fifo_store[4][12] ;
 wire \fifo0.fifo_store[4][13] ;
 wire \fifo0.fifo_store[4][14] ;
 wire \fifo0.fifo_store[4][15] ;
 wire \fifo0.fifo_store[4][1] ;
 wire \fifo0.fifo_store[4][2] ;
 wire \fifo0.fifo_store[4][3] ;
 wire \fifo0.fifo_store[4][4] ;
 wire \fifo0.fifo_store[4][5] ;
 wire \fifo0.fifo_store[4][6] ;
 wire \fifo0.fifo_store[4][7] ;
 wire \fifo0.fifo_store[4][8] ;
 wire \fifo0.fifo_store[4][9] ;
 wire \fifo0.fifo_store[50][0] ;
 wire \fifo0.fifo_store[50][10] ;
 wire \fifo0.fifo_store[50][11] ;
 wire \fifo0.fifo_store[50][12] ;
 wire \fifo0.fifo_store[50][13] ;
 wire \fifo0.fifo_store[50][14] ;
 wire \fifo0.fifo_store[50][15] ;
 wire \fifo0.fifo_store[50][1] ;
 wire \fifo0.fifo_store[50][2] ;
 wire \fifo0.fifo_store[50][3] ;
 wire \fifo0.fifo_store[50][4] ;
 wire \fifo0.fifo_store[50][5] ;
 wire \fifo0.fifo_store[50][6] ;
 wire \fifo0.fifo_store[50][7] ;
 wire \fifo0.fifo_store[50][8] ;
 wire \fifo0.fifo_store[50][9] ;
 wire \fifo0.fifo_store[51][0] ;
 wire \fifo0.fifo_store[51][10] ;
 wire \fifo0.fifo_store[51][11] ;
 wire \fifo0.fifo_store[51][12] ;
 wire \fifo0.fifo_store[51][13] ;
 wire \fifo0.fifo_store[51][14] ;
 wire \fifo0.fifo_store[51][15] ;
 wire \fifo0.fifo_store[51][1] ;
 wire \fifo0.fifo_store[51][2] ;
 wire \fifo0.fifo_store[51][3] ;
 wire \fifo0.fifo_store[51][4] ;
 wire \fifo0.fifo_store[51][5] ;
 wire \fifo0.fifo_store[51][6] ;
 wire \fifo0.fifo_store[51][7] ;
 wire \fifo0.fifo_store[51][8] ;
 wire \fifo0.fifo_store[51][9] ;
 wire \fifo0.fifo_store[52][0] ;
 wire \fifo0.fifo_store[52][10] ;
 wire \fifo0.fifo_store[52][11] ;
 wire \fifo0.fifo_store[52][12] ;
 wire \fifo0.fifo_store[52][13] ;
 wire \fifo0.fifo_store[52][14] ;
 wire \fifo0.fifo_store[52][15] ;
 wire \fifo0.fifo_store[52][1] ;
 wire \fifo0.fifo_store[52][2] ;
 wire \fifo0.fifo_store[52][3] ;
 wire \fifo0.fifo_store[52][4] ;
 wire \fifo0.fifo_store[52][5] ;
 wire \fifo0.fifo_store[52][6] ;
 wire \fifo0.fifo_store[52][7] ;
 wire \fifo0.fifo_store[52][8] ;
 wire \fifo0.fifo_store[52][9] ;
 wire \fifo0.fifo_store[53][0] ;
 wire \fifo0.fifo_store[53][10] ;
 wire \fifo0.fifo_store[53][11] ;
 wire \fifo0.fifo_store[53][12] ;
 wire \fifo0.fifo_store[53][13] ;
 wire \fifo0.fifo_store[53][14] ;
 wire \fifo0.fifo_store[53][15] ;
 wire \fifo0.fifo_store[53][1] ;
 wire \fifo0.fifo_store[53][2] ;
 wire \fifo0.fifo_store[53][3] ;
 wire \fifo0.fifo_store[53][4] ;
 wire \fifo0.fifo_store[53][5] ;
 wire \fifo0.fifo_store[53][6] ;
 wire \fifo0.fifo_store[53][7] ;
 wire \fifo0.fifo_store[53][8] ;
 wire \fifo0.fifo_store[53][9] ;
 wire \fifo0.fifo_store[54][0] ;
 wire \fifo0.fifo_store[54][10] ;
 wire \fifo0.fifo_store[54][11] ;
 wire \fifo0.fifo_store[54][12] ;
 wire \fifo0.fifo_store[54][13] ;
 wire \fifo0.fifo_store[54][14] ;
 wire \fifo0.fifo_store[54][15] ;
 wire \fifo0.fifo_store[54][1] ;
 wire \fifo0.fifo_store[54][2] ;
 wire \fifo0.fifo_store[54][3] ;
 wire \fifo0.fifo_store[54][4] ;
 wire \fifo0.fifo_store[54][5] ;
 wire \fifo0.fifo_store[54][6] ;
 wire \fifo0.fifo_store[54][7] ;
 wire \fifo0.fifo_store[54][8] ;
 wire \fifo0.fifo_store[54][9] ;
 wire \fifo0.fifo_store[55][0] ;
 wire \fifo0.fifo_store[55][10] ;
 wire \fifo0.fifo_store[55][11] ;
 wire \fifo0.fifo_store[55][12] ;
 wire \fifo0.fifo_store[55][13] ;
 wire \fifo0.fifo_store[55][14] ;
 wire \fifo0.fifo_store[55][15] ;
 wire \fifo0.fifo_store[55][1] ;
 wire \fifo0.fifo_store[55][2] ;
 wire \fifo0.fifo_store[55][3] ;
 wire \fifo0.fifo_store[55][4] ;
 wire \fifo0.fifo_store[55][5] ;
 wire \fifo0.fifo_store[55][6] ;
 wire \fifo0.fifo_store[55][7] ;
 wire \fifo0.fifo_store[55][8] ;
 wire \fifo0.fifo_store[55][9] ;
 wire \fifo0.fifo_store[56][0] ;
 wire \fifo0.fifo_store[56][10] ;
 wire \fifo0.fifo_store[56][11] ;
 wire \fifo0.fifo_store[56][12] ;
 wire \fifo0.fifo_store[56][13] ;
 wire \fifo0.fifo_store[56][14] ;
 wire \fifo0.fifo_store[56][15] ;
 wire \fifo0.fifo_store[56][1] ;
 wire \fifo0.fifo_store[56][2] ;
 wire \fifo0.fifo_store[56][3] ;
 wire \fifo0.fifo_store[56][4] ;
 wire \fifo0.fifo_store[56][5] ;
 wire \fifo0.fifo_store[56][6] ;
 wire \fifo0.fifo_store[56][7] ;
 wire \fifo0.fifo_store[56][8] ;
 wire \fifo0.fifo_store[56][9] ;
 wire \fifo0.fifo_store[57][0] ;
 wire \fifo0.fifo_store[57][10] ;
 wire \fifo0.fifo_store[57][11] ;
 wire \fifo0.fifo_store[57][12] ;
 wire \fifo0.fifo_store[57][13] ;
 wire \fifo0.fifo_store[57][14] ;
 wire \fifo0.fifo_store[57][15] ;
 wire \fifo0.fifo_store[57][1] ;
 wire \fifo0.fifo_store[57][2] ;
 wire \fifo0.fifo_store[57][3] ;
 wire \fifo0.fifo_store[57][4] ;
 wire \fifo0.fifo_store[57][5] ;
 wire \fifo0.fifo_store[57][6] ;
 wire \fifo0.fifo_store[57][7] ;
 wire \fifo0.fifo_store[57][8] ;
 wire \fifo0.fifo_store[57][9] ;
 wire \fifo0.fifo_store[58][0] ;
 wire \fifo0.fifo_store[58][10] ;
 wire \fifo0.fifo_store[58][11] ;
 wire \fifo0.fifo_store[58][12] ;
 wire \fifo0.fifo_store[58][13] ;
 wire \fifo0.fifo_store[58][14] ;
 wire \fifo0.fifo_store[58][15] ;
 wire \fifo0.fifo_store[58][1] ;
 wire \fifo0.fifo_store[58][2] ;
 wire \fifo0.fifo_store[58][3] ;
 wire \fifo0.fifo_store[58][4] ;
 wire \fifo0.fifo_store[58][5] ;
 wire \fifo0.fifo_store[58][6] ;
 wire \fifo0.fifo_store[58][7] ;
 wire \fifo0.fifo_store[58][8] ;
 wire \fifo0.fifo_store[58][9] ;
 wire \fifo0.fifo_store[59][0] ;
 wire \fifo0.fifo_store[59][10] ;
 wire \fifo0.fifo_store[59][11] ;
 wire \fifo0.fifo_store[59][12] ;
 wire \fifo0.fifo_store[59][13] ;
 wire \fifo0.fifo_store[59][14] ;
 wire \fifo0.fifo_store[59][15] ;
 wire \fifo0.fifo_store[59][1] ;
 wire \fifo0.fifo_store[59][2] ;
 wire \fifo0.fifo_store[59][3] ;
 wire \fifo0.fifo_store[59][4] ;
 wire \fifo0.fifo_store[59][5] ;
 wire \fifo0.fifo_store[59][6] ;
 wire \fifo0.fifo_store[59][7] ;
 wire \fifo0.fifo_store[59][8] ;
 wire \fifo0.fifo_store[59][9] ;
 wire \fifo0.fifo_store[5][0] ;
 wire \fifo0.fifo_store[5][10] ;
 wire \fifo0.fifo_store[5][11] ;
 wire \fifo0.fifo_store[5][12] ;
 wire \fifo0.fifo_store[5][13] ;
 wire \fifo0.fifo_store[5][14] ;
 wire \fifo0.fifo_store[5][15] ;
 wire \fifo0.fifo_store[5][1] ;
 wire \fifo0.fifo_store[5][2] ;
 wire \fifo0.fifo_store[5][3] ;
 wire \fifo0.fifo_store[5][4] ;
 wire \fifo0.fifo_store[5][5] ;
 wire \fifo0.fifo_store[5][6] ;
 wire \fifo0.fifo_store[5][7] ;
 wire \fifo0.fifo_store[5][8] ;
 wire \fifo0.fifo_store[5][9] ;
 wire \fifo0.fifo_store[60][0] ;
 wire \fifo0.fifo_store[60][10] ;
 wire \fifo0.fifo_store[60][11] ;
 wire \fifo0.fifo_store[60][12] ;
 wire \fifo0.fifo_store[60][13] ;
 wire \fifo0.fifo_store[60][14] ;
 wire \fifo0.fifo_store[60][15] ;
 wire \fifo0.fifo_store[60][1] ;
 wire \fifo0.fifo_store[60][2] ;
 wire \fifo0.fifo_store[60][3] ;
 wire \fifo0.fifo_store[60][4] ;
 wire \fifo0.fifo_store[60][5] ;
 wire \fifo0.fifo_store[60][6] ;
 wire \fifo0.fifo_store[60][7] ;
 wire \fifo0.fifo_store[60][8] ;
 wire \fifo0.fifo_store[60][9] ;
 wire \fifo0.fifo_store[61][0] ;
 wire \fifo0.fifo_store[61][10] ;
 wire \fifo0.fifo_store[61][11] ;
 wire \fifo0.fifo_store[61][12] ;
 wire \fifo0.fifo_store[61][13] ;
 wire \fifo0.fifo_store[61][14] ;
 wire \fifo0.fifo_store[61][15] ;
 wire \fifo0.fifo_store[61][1] ;
 wire \fifo0.fifo_store[61][2] ;
 wire \fifo0.fifo_store[61][3] ;
 wire \fifo0.fifo_store[61][4] ;
 wire \fifo0.fifo_store[61][5] ;
 wire \fifo0.fifo_store[61][6] ;
 wire \fifo0.fifo_store[61][7] ;
 wire \fifo0.fifo_store[61][8] ;
 wire \fifo0.fifo_store[61][9] ;
 wire \fifo0.fifo_store[62][0] ;
 wire \fifo0.fifo_store[62][10] ;
 wire \fifo0.fifo_store[62][11] ;
 wire \fifo0.fifo_store[62][12] ;
 wire \fifo0.fifo_store[62][13] ;
 wire \fifo0.fifo_store[62][14] ;
 wire \fifo0.fifo_store[62][15] ;
 wire \fifo0.fifo_store[62][1] ;
 wire \fifo0.fifo_store[62][2] ;
 wire \fifo0.fifo_store[62][3] ;
 wire \fifo0.fifo_store[62][4] ;
 wire \fifo0.fifo_store[62][5] ;
 wire \fifo0.fifo_store[62][6] ;
 wire \fifo0.fifo_store[62][7] ;
 wire \fifo0.fifo_store[62][8] ;
 wire \fifo0.fifo_store[62][9] ;
 wire \fifo0.fifo_store[63][0] ;
 wire \fifo0.fifo_store[63][10] ;
 wire \fifo0.fifo_store[63][11] ;
 wire \fifo0.fifo_store[63][12] ;
 wire \fifo0.fifo_store[63][13] ;
 wire \fifo0.fifo_store[63][14] ;
 wire \fifo0.fifo_store[63][15] ;
 wire \fifo0.fifo_store[63][1] ;
 wire \fifo0.fifo_store[63][2] ;
 wire \fifo0.fifo_store[63][3] ;
 wire \fifo0.fifo_store[63][4] ;
 wire \fifo0.fifo_store[63][5] ;
 wire \fifo0.fifo_store[63][6] ;
 wire \fifo0.fifo_store[63][7] ;
 wire \fifo0.fifo_store[63][8] ;
 wire \fifo0.fifo_store[63][9] ;
 wire \fifo0.fifo_store[64][0] ;
 wire \fifo0.fifo_store[64][10] ;
 wire \fifo0.fifo_store[64][11] ;
 wire \fifo0.fifo_store[64][12] ;
 wire \fifo0.fifo_store[64][13] ;
 wire \fifo0.fifo_store[64][14] ;
 wire \fifo0.fifo_store[64][15] ;
 wire \fifo0.fifo_store[64][1] ;
 wire \fifo0.fifo_store[64][2] ;
 wire \fifo0.fifo_store[64][3] ;
 wire \fifo0.fifo_store[64][4] ;
 wire \fifo0.fifo_store[64][5] ;
 wire \fifo0.fifo_store[64][6] ;
 wire \fifo0.fifo_store[64][7] ;
 wire \fifo0.fifo_store[64][8] ;
 wire \fifo0.fifo_store[64][9] ;
 wire \fifo0.fifo_store[65][0] ;
 wire \fifo0.fifo_store[65][10] ;
 wire \fifo0.fifo_store[65][11] ;
 wire \fifo0.fifo_store[65][12] ;
 wire \fifo0.fifo_store[65][13] ;
 wire \fifo0.fifo_store[65][14] ;
 wire \fifo0.fifo_store[65][15] ;
 wire \fifo0.fifo_store[65][1] ;
 wire \fifo0.fifo_store[65][2] ;
 wire \fifo0.fifo_store[65][3] ;
 wire \fifo0.fifo_store[65][4] ;
 wire \fifo0.fifo_store[65][5] ;
 wire \fifo0.fifo_store[65][6] ;
 wire \fifo0.fifo_store[65][7] ;
 wire \fifo0.fifo_store[65][8] ;
 wire \fifo0.fifo_store[65][9] ;
 wire \fifo0.fifo_store[66][0] ;
 wire \fifo0.fifo_store[66][10] ;
 wire \fifo0.fifo_store[66][11] ;
 wire \fifo0.fifo_store[66][12] ;
 wire \fifo0.fifo_store[66][13] ;
 wire \fifo0.fifo_store[66][14] ;
 wire \fifo0.fifo_store[66][15] ;
 wire \fifo0.fifo_store[66][1] ;
 wire \fifo0.fifo_store[66][2] ;
 wire \fifo0.fifo_store[66][3] ;
 wire \fifo0.fifo_store[66][4] ;
 wire \fifo0.fifo_store[66][5] ;
 wire \fifo0.fifo_store[66][6] ;
 wire \fifo0.fifo_store[66][7] ;
 wire \fifo0.fifo_store[66][8] ;
 wire \fifo0.fifo_store[66][9] ;
 wire \fifo0.fifo_store[67][0] ;
 wire \fifo0.fifo_store[67][10] ;
 wire \fifo0.fifo_store[67][11] ;
 wire \fifo0.fifo_store[67][12] ;
 wire \fifo0.fifo_store[67][13] ;
 wire \fifo0.fifo_store[67][14] ;
 wire \fifo0.fifo_store[67][15] ;
 wire \fifo0.fifo_store[67][1] ;
 wire \fifo0.fifo_store[67][2] ;
 wire \fifo0.fifo_store[67][3] ;
 wire \fifo0.fifo_store[67][4] ;
 wire \fifo0.fifo_store[67][5] ;
 wire \fifo0.fifo_store[67][6] ;
 wire \fifo0.fifo_store[67][7] ;
 wire \fifo0.fifo_store[67][8] ;
 wire \fifo0.fifo_store[67][9] ;
 wire \fifo0.fifo_store[68][0] ;
 wire \fifo0.fifo_store[68][10] ;
 wire \fifo0.fifo_store[68][11] ;
 wire \fifo0.fifo_store[68][12] ;
 wire \fifo0.fifo_store[68][13] ;
 wire \fifo0.fifo_store[68][14] ;
 wire \fifo0.fifo_store[68][15] ;
 wire \fifo0.fifo_store[68][1] ;
 wire \fifo0.fifo_store[68][2] ;
 wire \fifo0.fifo_store[68][3] ;
 wire \fifo0.fifo_store[68][4] ;
 wire \fifo0.fifo_store[68][5] ;
 wire \fifo0.fifo_store[68][6] ;
 wire \fifo0.fifo_store[68][7] ;
 wire \fifo0.fifo_store[68][8] ;
 wire \fifo0.fifo_store[68][9] ;
 wire \fifo0.fifo_store[69][0] ;
 wire \fifo0.fifo_store[69][10] ;
 wire \fifo0.fifo_store[69][11] ;
 wire \fifo0.fifo_store[69][12] ;
 wire \fifo0.fifo_store[69][13] ;
 wire \fifo0.fifo_store[69][14] ;
 wire \fifo0.fifo_store[69][15] ;
 wire \fifo0.fifo_store[69][1] ;
 wire \fifo0.fifo_store[69][2] ;
 wire \fifo0.fifo_store[69][3] ;
 wire \fifo0.fifo_store[69][4] ;
 wire \fifo0.fifo_store[69][5] ;
 wire \fifo0.fifo_store[69][6] ;
 wire \fifo0.fifo_store[69][7] ;
 wire \fifo0.fifo_store[69][8] ;
 wire \fifo0.fifo_store[69][9] ;
 wire \fifo0.fifo_store[6][0] ;
 wire \fifo0.fifo_store[6][10] ;
 wire \fifo0.fifo_store[6][11] ;
 wire \fifo0.fifo_store[6][12] ;
 wire \fifo0.fifo_store[6][13] ;
 wire \fifo0.fifo_store[6][14] ;
 wire \fifo0.fifo_store[6][15] ;
 wire \fifo0.fifo_store[6][1] ;
 wire \fifo0.fifo_store[6][2] ;
 wire \fifo0.fifo_store[6][3] ;
 wire \fifo0.fifo_store[6][4] ;
 wire \fifo0.fifo_store[6][5] ;
 wire \fifo0.fifo_store[6][6] ;
 wire \fifo0.fifo_store[6][7] ;
 wire \fifo0.fifo_store[6][8] ;
 wire \fifo0.fifo_store[6][9] ;
 wire \fifo0.fifo_store[70][0] ;
 wire \fifo0.fifo_store[70][10] ;
 wire \fifo0.fifo_store[70][11] ;
 wire \fifo0.fifo_store[70][12] ;
 wire \fifo0.fifo_store[70][13] ;
 wire \fifo0.fifo_store[70][14] ;
 wire \fifo0.fifo_store[70][15] ;
 wire \fifo0.fifo_store[70][1] ;
 wire \fifo0.fifo_store[70][2] ;
 wire \fifo0.fifo_store[70][3] ;
 wire \fifo0.fifo_store[70][4] ;
 wire \fifo0.fifo_store[70][5] ;
 wire \fifo0.fifo_store[70][6] ;
 wire \fifo0.fifo_store[70][7] ;
 wire \fifo0.fifo_store[70][8] ;
 wire \fifo0.fifo_store[70][9] ;
 wire \fifo0.fifo_store[71][0] ;
 wire \fifo0.fifo_store[71][10] ;
 wire \fifo0.fifo_store[71][11] ;
 wire \fifo0.fifo_store[71][12] ;
 wire \fifo0.fifo_store[71][13] ;
 wire \fifo0.fifo_store[71][14] ;
 wire \fifo0.fifo_store[71][15] ;
 wire \fifo0.fifo_store[71][1] ;
 wire \fifo0.fifo_store[71][2] ;
 wire \fifo0.fifo_store[71][3] ;
 wire \fifo0.fifo_store[71][4] ;
 wire \fifo0.fifo_store[71][5] ;
 wire \fifo0.fifo_store[71][6] ;
 wire \fifo0.fifo_store[71][7] ;
 wire \fifo0.fifo_store[71][8] ;
 wire \fifo0.fifo_store[71][9] ;
 wire \fifo0.fifo_store[72][0] ;
 wire \fifo0.fifo_store[72][10] ;
 wire \fifo0.fifo_store[72][11] ;
 wire \fifo0.fifo_store[72][12] ;
 wire \fifo0.fifo_store[72][13] ;
 wire \fifo0.fifo_store[72][14] ;
 wire \fifo0.fifo_store[72][15] ;
 wire \fifo0.fifo_store[72][1] ;
 wire \fifo0.fifo_store[72][2] ;
 wire \fifo0.fifo_store[72][3] ;
 wire \fifo0.fifo_store[72][4] ;
 wire \fifo0.fifo_store[72][5] ;
 wire \fifo0.fifo_store[72][6] ;
 wire \fifo0.fifo_store[72][7] ;
 wire \fifo0.fifo_store[72][8] ;
 wire \fifo0.fifo_store[72][9] ;
 wire \fifo0.fifo_store[73][0] ;
 wire \fifo0.fifo_store[73][10] ;
 wire \fifo0.fifo_store[73][11] ;
 wire \fifo0.fifo_store[73][12] ;
 wire \fifo0.fifo_store[73][13] ;
 wire \fifo0.fifo_store[73][14] ;
 wire \fifo0.fifo_store[73][15] ;
 wire \fifo0.fifo_store[73][1] ;
 wire \fifo0.fifo_store[73][2] ;
 wire \fifo0.fifo_store[73][3] ;
 wire \fifo0.fifo_store[73][4] ;
 wire \fifo0.fifo_store[73][5] ;
 wire \fifo0.fifo_store[73][6] ;
 wire \fifo0.fifo_store[73][7] ;
 wire \fifo0.fifo_store[73][8] ;
 wire \fifo0.fifo_store[73][9] ;
 wire \fifo0.fifo_store[74][0] ;
 wire \fifo0.fifo_store[74][10] ;
 wire \fifo0.fifo_store[74][11] ;
 wire \fifo0.fifo_store[74][12] ;
 wire \fifo0.fifo_store[74][13] ;
 wire \fifo0.fifo_store[74][14] ;
 wire \fifo0.fifo_store[74][15] ;
 wire \fifo0.fifo_store[74][1] ;
 wire \fifo0.fifo_store[74][2] ;
 wire \fifo0.fifo_store[74][3] ;
 wire \fifo0.fifo_store[74][4] ;
 wire \fifo0.fifo_store[74][5] ;
 wire \fifo0.fifo_store[74][6] ;
 wire \fifo0.fifo_store[74][7] ;
 wire \fifo0.fifo_store[74][8] ;
 wire \fifo0.fifo_store[74][9] ;
 wire \fifo0.fifo_store[75][0] ;
 wire \fifo0.fifo_store[75][10] ;
 wire \fifo0.fifo_store[75][11] ;
 wire \fifo0.fifo_store[75][12] ;
 wire \fifo0.fifo_store[75][13] ;
 wire \fifo0.fifo_store[75][14] ;
 wire \fifo0.fifo_store[75][15] ;
 wire \fifo0.fifo_store[75][1] ;
 wire \fifo0.fifo_store[75][2] ;
 wire \fifo0.fifo_store[75][3] ;
 wire \fifo0.fifo_store[75][4] ;
 wire \fifo0.fifo_store[75][5] ;
 wire \fifo0.fifo_store[75][6] ;
 wire \fifo0.fifo_store[75][7] ;
 wire \fifo0.fifo_store[75][8] ;
 wire \fifo0.fifo_store[75][9] ;
 wire \fifo0.fifo_store[76][0] ;
 wire \fifo0.fifo_store[76][10] ;
 wire \fifo0.fifo_store[76][11] ;
 wire \fifo0.fifo_store[76][12] ;
 wire \fifo0.fifo_store[76][13] ;
 wire \fifo0.fifo_store[76][14] ;
 wire \fifo0.fifo_store[76][15] ;
 wire \fifo0.fifo_store[76][1] ;
 wire \fifo0.fifo_store[76][2] ;
 wire \fifo0.fifo_store[76][3] ;
 wire \fifo0.fifo_store[76][4] ;
 wire \fifo0.fifo_store[76][5] ;
 wire \fifo0.fifo_store[76][6] ;
 wire \fifo0.fifo_store[76][7] ;
 wire \fifo0.fifo_store[76][8] ;
 wire \fifo0.fifo_store[76][9] ;
 wire \fifo0.fifo_store[77][0] ;
 wire \fifo0.fifo_store[77][10] ;
 wire \fifo0.fifo_store[77][11] ;
 wire \fifo0.fifo_store[77][12] ;
 wire \fifo0.fifo_store[77][13] ;
 wire \fifo0.fifo_store[77][14] ;
 wire \fifo0.fifo_store[77][15] ;
 wire \fifo0.fifo_store[77][1] ;
 wire \fifo0.fifo_store[77][2] ;
 wire \fifo0.fifo_store[77][3] ;
 wire \fifo0.fifo_store[77][4] ;
 wire \fifo0.fifo_store[77][5] ;
 wire \fifo0.fifo_store[77][6] ;
 wire \fifo0.fifo_store[77][7] ;
 wire \fifo0.fifo_store[77][8] ;
 wire \fifo0.fifo_store[77][9] ;
 wire \fifo0.fifo_store[78][0] ;
 wire \fifo0.fifo_store[78][10] ;
 wire \fifo0.fifo_store[78][11] ;
 wire \fifo0.fifo_store[78][12] ;
 wire \fifo0.fifo_store[78][13] ;
 wire \fifo0.fifo_store[78][14] ;
 wire \fifo0.fifo_store[78][15] ;
 wire \fifo0.fifo_store[78][1] ;
 wire \fifo0.fifo_store[78][2] ;
 wire \fifo0.fifo_store[78][3] ;
 wire \fifo0.fifo_store[78][4] ;
 wire \fifo0.fifo_store[78][5] ;
 wire \fifo0.fifo_store[78][6] ;
 wire \fifo0.fifo_store[78][7] ;
 wire \fifo0.fifo_store[78][8] ;
 wire \fifo0.fifo_store[78][9] ;
 wire \fifo0.fifo_store[79][0] ;
 wire \fifo0.fifo_store[79][10] ;
 wire \fifo0.fifo_store[79][11] ;
 wire \fifo0.fifo_store[79][12] ;
 wire \fifo0.fifo_store[79][13] ;
 wire \fifo0.fifo_store[79][14] ;
 wire \fifo0.fifo_store[79][15] ;
 wire \fifo0.fifo_store[79][1] ;
 wire \fifo0.fifo_store[79][2] ;
 wire \fifo0.fifo_store[79][3] ;
 wire \fifo0.fifo_store[79][4] ;
 wire \fifo0.fifo_store[79][5] ;
 wire \fifo0.fifo_store[79][6] ;
 wire \fifo0.fifo_store[79][7] ;
 wire \fifo0.fifo_store[79][8] ;
 wire \fifo0.fifo_store[79][9] ;
 wire \fifo0.fifo_store[7][0] ;
 wire \fifo0.fifo_store[7][10] ;
 wire \fifo0.fifo_store[7][11] ;
 wire \fifo0.fifo_store[7][12] ;
 wire \fifo0.fifo_store[7][13] ;
 wire \fifo0.fifo_store[7][14] ;
 wire \fifo0.fifo_store[7][15] ;
 wire \fifo0.fifo_store[7][1] ;
 wire \fifo0.fifo_store[7][2] ;
 wire \fifo0.fifo_store[7][3] ;
 wire \fifo0.fifo_store[7][4] ;
 wire \fifo0.fifo_store[7][5] ;
 wire \fifo0.fifo_store[7][6] ;
 wire \fifo0.fifo_store[7][7] ;
 wire \fifo0.fifo_store[7][8] ;
 wire \fifo0.fifo_store[7][9] ;
 wire \fifo0.fifo_store[80][0] ;
 wire \fifo0.fifo_store[80][10] ;
 wire \fifo0.fifo_store[80][11] ;
 wire \fifo0.fifo_store[80][12] ;
 wire \fifo0.fifo_store[80][13] ;
 wire \fifo0.fifo_store[80][14] ;
 wire \fifo0.fifo_store[80][15] ;
 wire \fifo0.fifo_store[80][1] ;
 wire \fifo0.fifo_store[80][2] ;
 wire \fifo0.fifo_store[80][3] ;
 wire \fifo0.fifo_store[80][4] ;
 wire \fifo0.fifo_store[80][5] ;
 wire \fifo0.fifo_store[80][6] ;
 wire \fifo0.fifo_store[80][7] ;
 wire \fifo0.fifo_store[80][8] ;
 wire \fifo0.fifo_store[80][9] ;
 wire \fifo0.fifo_store[81][0] ;
 wire \fifo0.fifo_store[81][10] ;
 wire \fifo0.fifo_store[81][11] ;
 wire \fifo0.fifo_store[81][12] ;
 wire \fifo0.fifo_store[81][13] ;
 wire \fifo0.fifo_store[81][14] ;
 wire \fifo0.fifo_store[81][15] ;
 wire \fifo0.fifo_store[81][1] ;
 wire \fifo0.fifo_store[81][2] ;
 wire \fifo0.fifo_store[81][3] ;
 wire \fifo0.fifo_store[81][4] ;
 wire \fifo0.fifo_store[81][5] ;
 wire \fifo0.fifo_store[81][6] ;
 wire \fifo0.fifo_store[81][7] ;
 wire \fifo0.fifo_store[81][8] ;
 wire \fifo0.fifo_store[81][9] ;
 wire \fifo0.fifo_store[82][0] ;
 wire \fifo0.fifo_store[82][10] ;
 wire \fifo0.fifo_store[82][11] ;
 wire \fifo0.fifo_store[82][12] ;
 wire \fifo0.fifo_store[82][13] ;
 wire \fifo0.fifo_store[82][14] ;
 wire \fifo0.fifo_store[82][15] ;
 wire \fifo0.fifo_store[82][1] ;
 wire \fifo0.fifo_store[82][2] ;
 wire \fifo0.fifo_store[82][3] ;
 wire \fifo0.fifo_store[82][4] ;
 wire \fifo0.fifo_store[82][5] ;
 wire \fifo0.fifo_store[82][6] ;
 wire \fifo0.fifo_store[82][7] ;
 wire \fifo0.fifo_store[82][8] ;
 wire \fifo0.fifo_store[82][9] ;
 wire \fifo0.fifo_store[83][0] ;
 wire \fifo0.fifo_store[83][10] ;
 wire \fifo0.fifo_store[83][11] ;
 wire \fifo0.fifo_store[83][12] ;
 wire \fifo0.fifo_store[83][13] ;
 wire \fifo0.fifo_store[83][14] ;
 wire \fifo0.fifo_store[83][15] ;
 wire \fifo0.fifo_store[83][1] ;
 wire \fifo0.fifo_store[83][2] ;
 wire \fifo0.fifo_store[83][3] ;
 wire \fifo0.fifo_store[83][4] ;
 wire \fifo0.fifo_store[83][5] ;
 wire \fifo0.fifo_store[83][6] ;
 wire \fifo0.fifo_store[83][7] ;
 wire \fifo0.fifo_store[83][8] ;
 wire \fifo0.fifo_store[83][9] ;
 wire \fifo0.fifo_store[84][0] ;
 wire \fifo0.fifo_store[84][10] ;
 wire \fifo0.fifo_store[84][11] ;
 wire \fifo0.fifo_store[84][12] ;
 wire \fifo0.fifo_store[84][13] ;
 wire \fifo0.fifo_store[84][14] ;
 wire \fifo0.fifo_store[84][15] ;
 wire \fifo0.fifo_store[84][1] ;
 wire \fifo0.fifo_store[84][2] ;
 wire \fifo0.fifo_store[84][3] ;
 wire \fifo0.fifo_store[84][4] ;
 wire \fifo0.fifo_store[84][5] ;
 wire \fifo0.fifo_store[84][6] ;
 wire \fifo0.fifo_store[84][7] ;
 wire \fifo0.fifo_store[84][8] ;
 wire \fifo0.fifo_store[84][9] ;
 wire \fifo0.fifo_store[85][0] ;
 wire \fifo0.fifo_store[85][10] ;
 wire \fifo0.fifo_store[85][11] ;
 wire \fifo0.fifo_store[85][12] ;
 wire \fifo0.fifo_store[85][13] ;
 wire \fifo0.fifo_store[85][14] ;
 wire \fifo0.fifo_store[85][15] ;
 wire \fifo0.fifo_store[85][1] ;
 wire \fifo0.fifo_store[85][2] ;
 wire \fifo0.fifo_store[85][3] ;
 wire \fifo0.fifo_store[85][4] ;
 wire \fifo0.fifo_store[85][5] ;
 wire \fifo0.fifo_store[85][6] ;
 wire \fifo0.fifo_store[85][7] ;
 wire \fifo0.fifo_store[85][8] ;
 wire \fifo0.fifo_store[85][9] ;
 wire \fifo0.fifo_store[86][0] ;
 wire \fifo0.fifo_store[86][10] ;
 wire \fifo0.fifo_store[86][11] ;
 wire \fifo0.fifo_store[86][12] ;
 wire \fifo0.fifo_store[86][13] ;
 wire \fifo0.fifo_store[86][14] ;
 wire \fifo0.fifo_store[86][15] ;
 wire \fifo0.fifo_store[86][1] ;
 wire \fifo0.fifo_store[86][2] ;
 wire \fifo0.fifo_store[86][3] ;
 wire \fifo0.fifo_store[86][4] ;
 wire \fifo0.fifo_store[86][5] ;
 wire \fifo0.fifo_store[86][6] ;
 wire \fifo0.fifo_store[86][7] ;
 wire \fifo0.fifo_store[86][8] ;
 wire \fifo0.fifo_store[86][9] ;
 wire \fifo0.fifo_store[87][0] ;
 wire \fifo0.fifo_store[87][10] ;
 wire \fifo0.fifo_store[87][11] ;
 wire \fifo0.fifo_store[87][12] ;
 wire \fifo0.fifo_store[87][13] ;
 wire \fifo0.fifo_store[87][14] ;
 wire \fifo0.fifo_store[87][15] ;
 wire \fifo0.fifo_store[87][1] ;
 wire \fifo0.fifo_store[87][2] ;
 wire \fifo0.fifo_store[87][3] ;
 wire \fifo0.fifo_store[87][4] ;
 wire \fifo0.fifo_store[87][5] ;
 wire \fifo0.fifo_store[87][6] ;
 wire \fifo0.fifo_store[87][7] ;
 wire \fifo0.fifo_store[87][8] ;
 wire \fifo0.fifo_store[87][9] ;
 wire \fifo0.fifo_store[88][0] ;
 wire \fifo0.fifo_store[88][10] ;
 wire \fifo0.fifo_store[88][11] ;
 wire \fifo0.fifo_store[88][12] ;
 wire \fifo0.fifo_store[88][13] ;
 wire \fifo0.fifo_store[88][14] ;
 wire \fifo0.fifo_store[88][15] ;
 wire \fifo0.fifo_store[88][1] ;
 wire \fifo0.fifo_store[88][2] ;
 wire \fifo0.fifo_store[88][3] ;
 wire \fifo0.fifo_store[88][4] ;
 wire \fifo0.fifo_store[88][5] ;
 wire \fifo0.fifo_store[88][6] ;
 wire \fifo0.fifo_store[88][7] ;
 wire \fifo0.fifo_store[88][8] ;
 wire \fifo0.fifo_store[88][9] ;
 wire \fifo0.fifo_store[89][0] ;
 wire \fifo0.fifo_store[89][10] ;
 wire \fifo0.fifo_store[89][11] ;
 wire \fifo0.fifo_store[89][12] ;
 wire \fifo0.fifo_store[89][13] ;
 wire \fifo0.fifo_store[89][14] ;
 wire \fifo0.fifo_store[89][15] ;
 wire \fifo0.fifo_store[89][1] ;
 wire \fifo0.fifo_store[89][2] ;
 wire \fifo0.fifo_store[89][3] ;
 wire \fifo0.fifo_store[89][4] ;
 wire \fifo0.fifo_store[89][5] ;
 wire \fifo0.fifo_store[89][6] ;
 wire \fifo0.fifo_store[89][7] ;
 wire \fifo0.fifo_store[89][8] ;
 wire \fifo0.fifo_store[89][9] ;
 wire \fifo0.fifo_store[8][0] ;
 wire \fifo0.fifo_store[8][10] ;
 wire \fifo0.fifo_store[8][11] ;
 wire \fifo0.fifo_store[8][12] ;
 wire \fifo0.fifo_store[8][13] ;
 wire \fifo0.fifo_store[8][14] ;
 wire \fifo0.fifo_store[8][15] ;
 wire \fifo0.fifo_store[8][1] ;
 wire \fifo0.fifo_store[8][2] ;
 wire \fifo0.fifo_store[8][3] ;
 wire \fifo0.fifo_store[8][4] ;
 wire \fifo0.fifo_store[8][5] ;
 wire \fifo0.fifo_store[8][6] ;
 wire \fifo0.fifo_store[8][7] ;
 wire \fifo0.fifo_store[8][8] ;
 wire \fifo0.fifo_store[8][9] ;
 wire \fifo0.fifo_store[90][0] ;
 wire \fifo0.fifo_store[90][10] ;
 wire \fifo0.fifo_store[90][11] ;
 wire \fifo0.fifo_store[90][12] ;
 wire \fifo0.fifo_store[90][13] ;
 wire \fifo0.fifo_store[90][14] ;
 wire \fifo0.fifo_store[90][15] ;
 wire \fifo0.fifo_store[90][1] ;
 wire \fifo0.fifo_store[90][2] ;
 wire \fifo0.fifo_store[90][3] ;
 wire \fifo0.fifo_store[90][4] ;
 wire \fifo0.fifo_store[90][5] ;
 wire \fifo0.fifo_store[90][6] ;
 wire \fifo0.fifo_store[90][7] ;
 wire \fifo0.fifo_store[90][8] ;
 wire \fifo0.fifo_store[90][9] ;
 wire \fifo0.fifo_store[91][0] ;
 wire \fifo0.fifo_store[91][10] ;
 wire \fifo0.fifo_store[91][11] ;
 wire \fifo0.fifo_store[91][12] ;
 wire \fifo0.fifo_store[91][13] ;
 wire \fifo0.fifo_store[91][14] ;
 wire \fifo0.fifo_store[91][15] ;
 wire \fifo0.fifo_store[91][1] ;
 wire \fifo0.fifo_store[91][2] ;
 wire \fifo0.fifo_store[91][3] ;
 wire \fifo0.fifo_store[91][4] ;
 wire \fifo0.fifo_store[91][5] ;
 wire \fifo0.fifo_store[91][6] ;
 wire \fifo0.fifo_store[91][7] ;
 wire \fifo0.fifo_store[91][8] ;
 wire \fifo0.fifo_store[91][9] ;
 wire \fifo0.fifo_store[92][0] ;
 wire \fifo0.fifo_store[92][10] ;
 wire \fifo0.fifo_store[92][11] ;
 wire \fifo0.fifo_store[92][12] ;
 wire \fifo0.fifo_store[92][13] ;
 wire \fifo0.fifo_store[92][14] ;
 wire \fifo0.fifo_store[92][15] ;
 wire \fifo0.fifo_store[92][1] ;
 wire \fifo0.fifo_store[92][2] ;
 wire \fifo0.fifo_store[92][3] ;
 wire \fifo0.fifo_store[92][4] ;
 wire \fifo0.fifo_store[92][5] ;
 wire \fifo0.fifo_store[92][6] ;
 wire \fifo0.fifo_store[92][7] ;
 wire \fifo0.fifo_store[92][8] ;
 wire \fifo0.fifo_store[92][9] ;
 wire \fifo0.fifo_store[93][0] ;
 wire \fifo0.fifo_store[93][10] ;
 wire \fifo0.fifo_store[93][11] ;
 wire \fifo0.fifo_store[93][12] ;
 wire \fifo0.fifo_store[93][13] ;
 wire \fifo0.fifo_store[93][14] ;
 wire \fifo0.fifo_store[93][15] ;
 wire \fifo0.fifo_store[93][1] ;
 wire \fifo0.fifo_store[93][2] ;
 wire \fifo0.fifo_store[93][3] ;
 wire \fifo0.fifo_store[93][4] ;
 wire \fifo0.fifo_store[93][5] ;
 wire \fifo0.fifo_store[93][6] ;
 wire \fifo0.fifo_store[93][7] ;
 wire \fifo0.fifo_store[93][8] ;
 wire \fifo0.fifo_store[93][9] ;
 wire \fifo0.fifo_store[94][0] ;
 wire \fifo0.fifo_store[94][10] ;
 wire \fifo0.fifo_store[94][11] ;
 wire \fifo0.fifo_store[94][12] ;
 wire \fifo0.fifo_store[94][13] ;
 wire \fifo0.fifo_store[94][14] ;
 wire \fifo0.fifo_store[94][15] ;
 wire \fifo0.fifo_store[94][1] ;
 wire \fifo0.fifo_store[94][2] ;
 wire \fifo0.fifo_store[94][3] ;
 wire \fifo0.fifo_store[94][4] ;
 wire \fifo0.fifo_store[94][5] ;
 wire \fifo0.fifo_store[94][6] ;
 wire \fifo0.fifo_store[94][7] ;
 wire \fifo0.fifo_store[94][8] ;
 wire \fifo0.fifo_store[94][9] ;
 wire \fifo0.fifo_store[95][0] ;
 wire \fifo0.fifo_store[95][10] ;
 wire \fifo0.fifo_store[95][11] ;
 wire \fifo0.fifo_store[95][12] ;
 wire \fifo0.fifo_store[95][13] ;
 wire \fifo0.fifo_store[95][14] ;
 wire \fifo0.fifo_store[95][15] ;
 wire \fifo0.fifo_store[95][1] ;
 wire \fifo0.fifo_store[95][2] ;
 wire \fifo0.fifo_store[95][3] ;
 wire \fifo0.fifo_store[95][4] ;
 wire \fifo0.fifo_store[95][5] ;
 wire \fifo0.fifo_store[95][6] ;
 wire \fifo0.fifo_store[95][7] ;
 wire \fifo0.fifo_store[95][8] ;
 wire \fifo0.fifo_store[95][9] ;
 wire \fifo0.fifo_store[96][0] ;
 wire \fifo0.fifo_store[96][10] ;
 wire \fifo0.fifo_store[96][11] ;
 wire \fifo0.fifo_store[96][12] ;
 wire \fifo0.fifo_store[96][13] ;
 wire \fifo0.fifo_store[96][14] ;
 wire \fifo0.fifo_store[96][15] ;
 wire \fifo0.fifo_store[96][1] ;
 wire \fifo0.fifo_store[96][2] ;
 wire \fifo0.fifo_store[96][3] ;
 wire \fifo0.fifo_store[96][4] ;
 wire \fifo0.fifo_store[96][5] ;
 wire \fifo0.fifo_store[96][6] ;
 wire \fifo0.fifo_store[96][7] ;
 wire \fifo0.fifo_store[96][8] ;
 wire \fifo0.fifo_store[96][9] ;
 wire \fifo0.fifo_store[97][0] ;
 wire \fifo0.fifo_store[97][10] ;
 wire \fifo0.fifo_store[97][11] ;
 wire \fifo0.fifo_store[97][12] ;
 wire \fifo0.fifo_store[97][13] ;
 wire \fifo0.fifo_store[97][14] ;
 wire \fifo0.fifo_store[97][15] ;
 wire \fifo0.fifo_store[97][1] ;
 wire \fifo0.fifo_store[97][2] ;
 wire \fifo0.fifo_store[97][3] ;
 wire \fifo0.fifo_store[97][4] ;
 wire \fifo0.fifo_store[97][5] ;
 wire \fifo0.fifo_store[97][6] ;
 wire \fifo0.fifo_store[97][7] ;
 wire \fifo0.fifo_store[97][8] ;
 wire \fifo0.fifo_store[97][9] ;
 wire \fifo0.fifo_store[98][0] ;
 wire \fifo0.fifo_store[98][10] ;
 wire \fifo0.fifo_store[98][11] ;
 wire \fifo0.fifo_store[98][12] ;
 wire \fifo0.fifo_store[98][13] ;
 wire \fifo0.fifo_store[98][14] ;
 wire \fifo0.fifo_store[98][15] ;
 wire \fifo0.fifo_store[98][1] ;
 wire \fifo0.fifo_store[98][2] ;
 wire \fifo0.fifo_store[98][3] ;
 wire \fifo0.fifo_store[98][4] ;
 wire \fifo0.fifo_store[98][5] ;
 wire \fifo0.fifo_store[98][6] ;
 wire \fifo0.fifo_store[98][7] ;
 wire \fifo0.fifo_store[98][8] ;
 wire \fifo0.fifo_store[98][9] ;
 wire \fifo0.fifo_store[99][0] ;
 wire \fifo0.fifo_store[99][10] ;
 wire \fifo0.fifo_store[99][11] ;
 wire \fifo0.fifo_store[99][12] ;
 wire \fifo0.fifo_store[99][13] ;
 wire \fifo0.fifo_store[99][14] ;
 wire \fifo0.fifo_store[99][15] ;
 wire \fifo0.fifo_store[99][1] ;
 wire \fifo0.fifo_store[99][2] ;
 wire \fifo0.fifo_store[99][3] ;
 wire \fifo0.fifo_store[99][4] ;
 wire \fifo0.fifo_store[99][5] ;
 wire \fifo0.fifo_store[99][6] ;
 wire \fifo0.fifo_store[99][7] ;
 wire \fifo0.fifo_store[99][8] ;
 wire \fifo0.fifo_store[99][9] ;
 wire \fifo0.fifo_store[9][0] ;
 wire \fifo0.fifo_store[9][10] ;
 wire \fifo0.fifo_store[9][11] ;
 wire \fifo0.fifo_store[9][12] ;
 wire \fifo0.fifo_store[9][13] ;
 wire \fifo0.fifo_store[9][14] ;
 wire \fifo0.fifo_store[9][15] ;
 wire \fifo0.fifo_store[9][1] ;
 wire \fifo0.fifo_store[9][2] ;
 wire \fifo0.fifo_store[9][3] ;
 wire \fifo0.fifo_store[9][4] ;
 wire \fifo0.fifo_store[9][5] ;
 wire \fifo0.fifo_store[9][6] ;
 wire \fifo0.fifo_store[9][7] ;
 wire \fifo0.fifo_store[9][8] ;
 wire \fifo0.fifo_store[9][9] ;
 wire \fifo0.read_ptr[0] ;
 wire \fifo0.read_ptr[1] ;
 wire \fifo0.read_ptr[2] ;
 wire \fifo0.read_ptr[3] ;
 wire \fifo0.read_ptr[4] ;
 wire \fifo0.read_ptr[5] ;
 wire \fifo0.read_ptr[6] ;
 wire \fifo0.write_ptr[0] ;
 wire \fifo0.write_ptr[1] ;
 wire \fifo0.write_ptr[2] ;
 wire \fifo0.write_ptr[3] ;
 wire \fifo0.write_ptr[4] ;
 wire \fifo0.write_ptr[5] ;
 wire \fifo0.write_ptr[6] ;
 wire \sinegen0.read_ptr[0] ;
 wire \sinegen0.read_ptr[1] ;
 wire \sinegen0.read_ptr[2] ;
 wire \sinegen0.read_ptr[3] ;
 wire \sinegen0.read_ptr[4] ;
 wire \sinegen0.read_ptr[5] ;
 wire \sinegen0.read_ptr[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_leaf_108_clk_i;
 wire clknet_leaf_109_clk_i;
 wire clknet_leaf_110_clk_i;
 wire clknet_leaf_111_clk_i;
 wire clknet_leaf_112_clk_i;
 wire clknet_leaf_113_clk_i;
 wire clknet_leaf_114_clk_i;
 wire clknet_leaf_115_clk_i;
 wire clknet_leaf_116_clk_i;
 wire clknet_leaf_117_clk_i;
 wire clknet_leaf_118_clk_i;
 wire clknet_leaf_119_clk_i;
 wire clknet_leaf_120_clk_i;
 wire clknet_leaf_121_clk_i;
 wire clknet_leaf_122_clk_i;
 wire clknet_leaf_123_clk_i;
 wire clknet_leaf_124_clk_i;
 wire clknet_leaf_125_clk_i;
 wire clknet_leaf_126_clk_i;
 wire clknet_leaf_127_clk_i;
 wire clknet_leaf_128_clk_i;
 wire clknet_leaf_129_clk_i;
 wire clknet_leaf_130_clk_i;
 wire clknet_leaf_131_clk_i;
 wire clknet_leaf_132_clk_i;
 wire clknet_leaf_133_clk_i;
 wire clknet_leaf_134_clk_i;
 wire clknet_leaf_135_clk_i;
 wire clknet_leaf_136_clk_i;
 wire clknet_leaf_137_clk_i;
 wire clknet_leaf_138_clk_i;
 wire clknet_leaf_139_clk_i;
 wire clknet_leaf_140_clk_i;
 wire clknet_leaf_141_clk_i;
 wire clknet_leaf_142_clk_i;
 wire clknet_leaf_143_clk_i;
 wire clknet_leaf_144_clk_i;
 wire clknet_leaf_145_clk_i;
 wire clknet_leaf_146_clk_i;
 wire clknet_leaf_147_clk_i;
 wire clknet_leaf_148_clk_i;
 wire clknet_leaf_149_clk_i;
 wire clknet_leaf_150_clk_i;
 wire clknet_leaf_151_clk_i;
 wire clknet_leaf_152_clk_i;
 wire clknet_leaf_153_clk_i;
 wire clknet_leaf_154_clk_i;
 wire clknet_leaf_155_clk_i;
 wire clknet_leaf_156_clk_i;
 wire clknet_leaf_157_clk_i;
 wire clknet_leaf_158_clk_i;
 wire clknet_leaf_159_clk_i;
 wire clknet_leaf_160_clk_i;
 wire clknet_leaf_161_clk_i;
 wire clknet_leaf_162_clk_i;
 wire clknet_leaf_163_clk_i;
 wire clknet_leaf_164_clk_i;
 wire clknet_leaf_165_clk_i;
 wire clknet_leaf_166_clk_i;
 wire clknet_leaf_167_clk_i;
 wire clknet_leaf_168_clk_i;
 wire clknet_leaf_169_clk_i;
 wire clknet_leaf_170_clk_i;
 wire clknet_leaf_171_clk_i;
 wire clknet_leaf_172_clk_i;
 wire clknet_leaf_173_clk_i;
 wire clknet_leaf_174_clk_i;
 wire clknet_leaf_175_clk_i;
 wire clknet_leaf_176_clk_i;
 wire clknet_leaf_177_clk_i;
 wire clknet_leaf_178_clk_i;
 wire clknet_leaf_179_clk_i;
 wire clknet_leaf_180_clk_i;
 wire clknet_leaf_181_clk_i;
 wire clknet_leaf_182_clk_i;
 wire clknet_leaf_183_clk_i;
 wire clknet_leaf_184_clk_i;
 wire clknet_leaf_185_clk_i;
 wire clknet_leaf_186_clk_i;
 wire clknet_leaf_187_clk_i;
 wire clknet_leaf_188_clk_i;
 wire clknet_leaf_189_clk_i;
 wire clknet_leaf_190_clk_i;
 wire clknet_leaf_191_clk_i;
 wire clknet_leaf_192_clk_i;
 wire clknet_leaf_193_clk_i;
 wire clknet_leaf_194_clk_i;
 wire clknet_leaf_195_clk_i;
 wire clknet_leaf_196_clk_i;
 wire clknet_leaf_197_clk_i;
 wire clknet_leaf_198_clk_i;
 wire clknet_leaf_199_clk_i;
 wire clknet_leaf_200_clk_i;
 wire clknet_leaf_201_clk_i;
 wire clknet_leaf_202_clk_i;
 wire clknet_leaf_203_clk_i;
 wire clknet_leaf_204_clk_i;
 wire clknet_leaf_205_clk_i;
 wire clknet_leaf_206_clk_i;
 wire clknet_leaf_207_clk_i;
 wire clknet_leaf_208_clk_i;
 wire clknet_leaf_209_clk_i;
 wire clknet_leaf_210_clk_i;
 wire clknet_leaf_211_clk_i;
 wire clknet_leaf_212_clk_i;
 wire clknet_leaf_213_clk_i;
 wire clknet_leaf_214_clk_i;
 wire clknet_leaf_215_clk_i;
 wire clknet_leaf_216_clk_i;
 wire clknet_leaf_217_clk_i;
 wire clknet_leaf_218_clk_i;
 wire clknet_leaf_219_clk_i;
 wire clknet_leaf_220_clk_i;
 wire clknet_leaf_221_clk_i;
 wire clknet_leaf_222_clk_i;
 wire clknet_leaf_223_clk_i;
 wire clknet_leaf_224_clk_i;
 wire clknet_leaf_225_clk_i;
 wire clknet_leaf_226_clk_i;
 wire clknet_leaf_227_clk_i;
 wire clknet_leaf_228_clk_i;
 wire clknet_leaf_229_clk_i;
 wire clknet_leaf_230_clk_i;
 wire clknet_leaf_231_clk_i;
 wire clknet_leaf_232_clk_i;
 wire clknet_leaf_233_clk_i;
 wire clknet_leaf_234_clk_i;
 wire clknet_leaf_235_clk_i;
 wire clknet_leaf_236_clk_i;
 wire clknet_leaf_237_clk_i;
 wire clknet_leaf_238_clk_i;
 wire clknet_leaf_239_clk_i;
 wire clknet_leaf_240_clk_i;
 wire clknet_leaf_241_clk_i;
 wire clknet_leaf_242_clk_i;
 wire clknet_leaf_243_clk_i;
 wire clknet_leaf_244_clk_i;
 wire clknet_leaf_245_clk_i;
 wire clknet_leaf_246_clk_i;
 wire clknet_leaf_247_clk_i;
 wire clknet_leaf_248_clk_i;
 wire clknet_leaf_249_clk_i;
 wire clknet_leaf_250_clk_i;
 wire clknet_leaf_251_clk_i;
 wire clknet_leaf_252_clk_i;
 wire clknet_leaf_253_clk_i;
 wire clknet_leaf_254_clk_i;
 wire clknet_leaf_255_clk_i;
 wire clknet_leaf_256_clk_i;
 wire clknet_leaf_257_clk_i;
 wire clknet_leaf_258_clk_i;
 wire clknet_leaf_259_clk_i;
 wire clknet_leaf_260_clk_i;
 wire clknet_leaf_261_clk_i;
 wire clknet_leaf_262_clk_i;
 wire clknet_leaf_263_clk_i;
 wire clknet_leaf_264_clk_i;
 wire clknet_leaf_265_clk_i;
 wire clknet_leaf_266_clk_i;
 wire clknet_leaf_267_clk_i;
 wire clknet_leaf_268_clk_i;
 wire clknet_leaf_269_clk_i;
 wire clknet_leaf_270_clk_i;
 wire clknet_leaf_271_clk_i;
 wire clknet_leaf_272_clk_i;
 wire clknet_leaf_273_clk_i;
 wire clknet_leaf_274_clk_i;
 wire clknet_leaf_275_clk_i;
 wire clknet_leaf_277_clk_i;
 wire clknet_leaf_278_clk_i;
 wire clknet_leaf_279_clk_i;
 wire clknet_leaf_280_clk_i;
 wire clknet_leaf_281_clk_i;
 wire clknet_leaf_282_clk_i;
 wire clknet_leaf_283_clk_i;
 wire clknet_leaf_284_clk_i;
 wire clknet_leaf_285_clk_i;
 wire clknet_leaf_286_clk_i;
 wire clknet_leaf_287_clk_i;
 wire clknet_leaf_288_clk_i;
 wire clknet_leaf_289_clk_i;
 wire clknet_leaf_290_clk_i;
 wire clknet_leaf_291_clk_i;
 wire clknet_leaf_292_clk_i;
 wire clknet_leaf_293_clk_i;
 wire clknet_leaf_294_clk_i;
 wire clknet_leaf_295_clk_i;
 wire clknet_leaf_296_clk_i;
 wire clknet_leaf_297_clk_i;
 wire clknet_leaf_298_clk_i;
 wire clknet_leaf_299_clk_i;
 wire clknet_leaf_300_clk_i;
 wire clknet_leaf_301_clk_i;
 wire clknet_leaf_302_clk_i;
 wire clknet_leaf_303_clk_i;
 wire clknet_leaf_304_clk_i;
 wire clknet_leaf_305_clk_i;
 wire clknet_leaf_306_clk_i;
 wire clknet_leaf_307_clk_i;
 wire clknet_leaf_308_clk_i;
 wire clknet_leaf_309_clk_i;
 wire clknet_leaf_310_clk_i;
 wire clknet_leaf_311_clk_i;
 wire clknet_leaf_312_clk_i;
 wire clknet_leaf_313_clk_i;
 wire clknet_leaf_314_clk_i;
 wire clknet_leaf_315_clk_i;
 wire clknet_leaf_316_clk_i;
 wire clknet_leaf_317_clk_i;
 wire clknet_leaf_318_clk_i;
 wire clknet_leaf_319_clk_i;
 wire clknet_leaf_320_clk_i;
 wire clknet_leaf_321_clk_i;
 wire clknet_leaf_322_clk_i;
 wire clknet_leaf_323_clk_i;
 wire clknet_leaf_324_clk_i;
 wire clknet_leaf_325_clk_i;
 wire clknet_leaf_326_clk_i;
 wire clknet_leaf_327_clk_i;
 wire clknet_leaf_328_clk_i;
 wire clknet_leaf_329_clk_i;
 wire clknet_leaf_330_clk_i;
 wire clknet_leaf_331_clk_i;
 wire clknet_leaf_332_clk_i;
 wire clknet_leaf_333_clk_i;
 wire clknet_leaf_335_clk_i;
 wire clknet_leaf_336_clk_i;
 wire clknet_leaf_337_clk_i;
 wire clknet_leaf_338_clk_i;
 wire clknet_leaf_339_clk_i;
 wire clknet_leaf_340_clk_i;
 wire clknet_leaf_341_clk_i;
 wire clknet_leaf_342_clk_i;
 wire clknet_leaf_343_clk_i;
 wire clknet_0_clk_i;
 wire clknet_1_0_0_clk_i;
 wire clknet_1_0_1_clk_i;
 wire clknet_1_1_0_clk_i;
 wire clknet_1_1_1_clk_i;
 wire clknet_2_0_0_clk_i;
 wire clknet_2_0_1_clk_i;
 wire clknet_2_1_0_clk_i;
 wire clknet_2_1_1_clk_i;
 wire clknet_2_2_0_clk_i;
 wire clknet_2_2_1_clk_i;
 wire clknet_2_3_0_clk_i;
 wire clknet_2_3_1_clk_i;
 wire clknet_3_0_0_clk_i;
 wire clknet_3_1_0_clk_i;
 wire clknet_3_2_0_clk_i;
 wire clknet_3_3_0_clk_i;
 wire clknet_3_4_0_clk_i;
 wire clknet_3_5_0_clk_i;
 wire clknet_3_6_0_clk_i;
 wire clknet_3_7_0_clk_i;
 wire clknet_4_0_0_clk_i;
 wire clknet_4_1_0_clk_i;
 wire clknet_4_2_0_clk_i;
 wire clknet_4_3_0_clk_i;
 wire clknet_4_4_0_clk_i;
 wire clknet_4_5_0_clk_i;
 wire clknet_4_6_0_clk_i;
 wire clknet_4_7_0_clk_i;
 wire clknet_4_8_0_clk_i;
 wire clknet_4_9_0_clk_i;
 wire clknet_4_10_0_clk_i;
 wire clknet_4_11_0_clk_i;
 wire clknet_4_12_0_clk_i;
 wire clknet_4_13_0_clk_i;
 wire clknet_4_14_0_clk_i;
 wire clknet_4_15_0_clk_i;
 wire clknet_5_0_0_clk_i;
 wire clknet_5_1_0_clk_i;
 wire clknet_5_2_0_clk_i;
 wire clknet_5_3_0_clk_i;
 wire clknet_5_4_0_clk_i;
 wire clknet_5_5_0_clk_i;
 wire clknet_5_6_0_clk_i;
 wire clknet_5_7_0_clk_i;
 wire clknet_5_8_0_clk_i;
 wire clknet_5_9_0_clk_i;
 wire clknet_5_10_0_clk_i;
 wire clknet_5_11_0_clk_i;
 wire clknet_5_12_0_clk_i;
 wire clknet_5_13_0_clk_i;
 wire clknet_5_14_0_clk_i;
 wire clknet_5_15_0_clk_i;
 wire clknet_5_16_0_clk_i;
 wire clknet_5_17_0_clk_i;
 wire clknet_5_18_0_clk_i;
 wire clknet_5_19_0_clk_i;
 wire clknet_5_20_0_clk_i;
 wire clknet_5_21_0_clk_i;
 wire clknet_5_22_0_clk_i;
 wire clknet_5_23_0_clk_i;
 wire clknet_5_24_0_clk_i;
 wire clknet_5_25_0_clk_i;
 wire clknet_5_26_0_clk_i;
 wire clknet_5_27_0_clk_i;
 wire clknet_5_28_0_clk_i;
 wire clknet_5_29_0_clk_i;
 wire clknet_5_30_0_clk_i;
 wire clknet_5_31_0_clk_i;

 sky130_fd_sc_hd__xor2_1 _07436_ (.A(\fifo0.read_ptr[1] ),
    .B(\fifo0.write_ptr[1] ),
    .X(_03771_));
 sky130_fd_sc_hd__xor2_1 _07437_ (.A(\fifo0.read_ptr[5] ),
    .B(\fifo0.write_ptr[5] ),
    .X(_03772_));
 sky130_fd_sc_hd__xor2_1 _07438_ (.A(\fifo0.read_ptr[6] ),
    .B(\fifo0.write_ptr[6] ),
    .X(_03773_));
 sky130_fd_sc_hd__xnor2_1 _07439_ (.A(\fifo0.read_ptr[3] ),
    .B(\fifo0.write_ptr[3] ),
    .Y(_03774_));
 sky130_fd_sc_hd__xnor2_1 _07440_ (.A(\fifo0.read_ptr[0] ),
    .B(\fifo0.write_ptr[0] ),
    .Y(_03775_));
 sky130_fd_sc_hd__xnor2_1 _07441_ (.A(\fifo0.read_ptr[4] ),
    .B(\fifo0.write_ptr[4] ),
    .Y(_03776_));
 sky130_fd_sc_hd__xnor2_1 _07442_ (.A(\fifo0.read_ptr[2] ),
    .B(\fifo0.write_ptr[2] ),
    .Y(_03777_));
 sky130_fd_sc_hd__and4_1 _07443_ (.A(_03774_),
    .B(_03775_),
    .C(_03776_),
    .D(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__or4b_4 _07444_ (.A(_03771_),
    .B(_03772_),
    .C(_03773_),
    .D_N(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__inv_2 _07445_ (.A(_03779_),
    .Y(net37));
 sky130_fd_sc_hd__and3_1 _07446_ (.A(\fifo0.write_ptr[2] ),
    .B(\fifo0.write_ptr[1] ),
    .C(\fifo0.write_ptr[0] ),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_4 _07447_ (.A(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__and3_1 _07448_ (.A(\fifo0.write_ptr[4] ),
    .B(\fifo0.write_ptr[3] ),
    .C(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__and2_1 _07449_ (.A(\fifo0.write_ptr[5] ),
    .B(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__xor2_1 _07450_ (.A(_03773_),
    .B(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__and2_1 _07451_ (.A(\fifo0.write_ptr[1] ),
    .B(\fifo0.write_ptr[0] ),
    .X(_03785_));
 sky130_fd_sc_hd__nor2_1 _07452_ (.A(\fifo0.write_ptr[1] ),
    .B(\fifo0.write_ptr[0] ),
    .Y(_03786_));
 sky130_fd_sc_hd__or2_1 _07453_ (.A(_03785_),
    .B(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(\fifo0.write_ptr[2] ),
    .B(_03785_),
    .Y(_03788_));
 sky130_fd_sc_hd__or2_1 _07455_ (.A(_03781_),
    .B(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__a221o_1 _07456_ (.A1(\fifo0.read_ptr[1] ),
    .A2(_03787_),
    .B1(_03789_),
    .B2(\fifo0.read_ptr[2] ),
    .C1(_03775_),
    .X(_03790_));
 sky130_fd_sc_hd__o22ai_1 _07457_ (.A1(_03774_),
    .A2(_03781_),
    .B1(_03787_),
    .B2(\fifo0.read_ptr[1] ),
    .Y(_03791_));
 sky130_fd_sc_hd__xor2_1 _07458_ (.A(_03772_),
    .B(_03782_),
    .X(_03792_));
 sky130_fd_sc_hd__a21oi_1 _07459_ (.A1(\fifo0.write_ptr[3] ),
    .A2(_03781_),
    .B1(\fifo0.write_ptr[4] ),
    .Y(_03793_));
 sky130_fd_sc_hd__or2_2 _07460_ (.A(_03782_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__xor2_1 _07461_ (.A(\fifo0.read_ptr[4] ),
    .B(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__o21ai_1 _07462_ (.A1(\fifo0.read_ptr[2] ),
    .A2(_03789_),
    .B1(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__a2111o_1 _07463_ (.A1(_03774_),
    .A2(_03781_),
    .B1(_03791_),
    .C1(_03792_),
    .D1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__or3_1 _07464_ (.A(_03784_),
    .B(_03790_),
    .C(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__inv_2 _07465_ (.A(_03798_),
    .Y(net38));
 sky130_fd_sc_hd__inv_2 _07466_ (.A(net35),
    .Y(net34));
 sky130_fd_sc_hd__inv_4 _07467_ (.A(net21),
    .Y(_03799_));
 sky130_fd_sc_hd__or3b_4 _07468_ (.A(net36),
    .B(net38),
    .C_N(\fifo0.fifo_rdy ),
    .X(_03800_));
 sky130_fd_sc_hd__or2_1 _07469_ (.A(_03799_),
    .B(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__clkbuf_4 _07470_ (.A(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _07471_ (.A(\fifo0.write_ptr[3] ),
    .B(_03781_),
    .Y(_03803_));
 sky130_fd_sc_hd__nor2_1 _07472_ (.A(_03802_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_03794_),
    .B(_03802_),
    .Y(_03805_));
 sky130_fd_sc_hd__or2_2 _07474_ (.A(_03804_),
    .B(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__nor2_1 _07475_ (.A(\fifo0.write_ptr[5] ),
    .B(_03782_),
    .Y(_03807_));
 sky130_fd_sc_hd__or2_1 _07476_ (.A(_03783_),
    .B(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__nor2_1 _07477_ (.A(_03802_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__xnor2_1 _07478_ (.A(\fifo0.write_ptr[6] ),
    .B(_03783_),
    .Y(_03810_));
 sky130_fd_sc_hd__nor2_1 _07479_ (.A(_03810_),
    .B(_03802_),
    .Y(_03811_));
 sky130_fd_sc_hd__or2_1 _07480_ (.A(_03809_),
    .B(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__or2_1 _07481_ (.A(_03806_),
    .B(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__buf_12 _07482_ (.A(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__nor2_8 _07483_ (.A(_03781_),
    .B(_03802_),
    .Y(_03815_));
 sky130_fd_sc_hd__buf_12 _07484_ (.A(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__nor2_8 _07485_ (.A(_03814_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__nor2_8 _07486_ (.A(_03799_),
    .B(_03800_),
    .Y(_03818_));
 sky130_fd_sc_hd__buf_8 _07487_ (.A(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _07488_ (.A(\fifo0.fifo_data[0] ),
    .B(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__buf_2 _07489_ (.A(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__buf_4 _07490_ (.A(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__and2_1 _07491_ (.A(net21),
    .B(_03800_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_4 _07492_ (.A(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__or3_1 _07493_ (.A(_03814_),
    .B(_03815_),
    .C(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_4 _07494_ (.A(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_4 _07495_ (.A(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__a22o_1 _07496_ (.A1(_03817_),
    .A2(_03822_),
    .B1(_03827_),
    .B2(\fifo0.fifo_store[0][0] ),
    .X(_00007_));
 sky130_fd_sc_hd__and2_1 _07497_ (.A(\fifo0.fifo_data[1] ),
    .B(_03818_),
    .X(_03828_));
 sky130_fd_sc_hd__buf_4 _07498_ (.A(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__buf_6 _07499_ (.A(_03817_),
    .X(_03830_));
 sky130_fd_sc_hd__a22o_1 _07500_ (.A1(\fifo0.fifo_store[0][1] ),
    .A2(_03827_),
    .B1(_03829_),
    .B2(_03830_),
    .X(_00008_));
 sky130_fd_sc_hd__and2_1 _07501_ (.A(\fifo0.fifo_data[2] ),
    .B(_03819_),
    .X(_03831_));
 sky130_fd_sc_hd__buf_4 _07502_ (.A(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__a22o_1 _07503_ (.A1(\fifo0.fifo_store[0][2] ),
    .A2(_03827_),
    .B1(_03832_),
    .B2(_03830_),
    .X(_00009_));
 sky130_fd_sc_hd__and2_1 _07504_ (.A(\fifo0.fifo_data[3] ),
    .B(_03819_),
    .X(_03833_));
 sky130_fd_sc_hd__buf_6 _07505_ (.A(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__a22o_1 _07506_ (.A1(\fifo0.fifo_store[0][3] ),
    .A2(_03827_),
    .B1(_03834_),
    .B2(_03830_),
    .X(_00010_));
 sky130_fd_sc_hd__and2_1 _07507_ (.A(\fifo0.fifo_data[4] ),
    .B(_03819_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_4 _07508_ (.A(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__a22o_1 _07509_ (.A1(\fifo0.fifo_store[0][4] ),
    .A2(_03827_),
    .B1(_03836_),
    .B2(_03830_),
    .X(_00011_));
 sky130_fd_sc_hd__and2_2 _07510_ (.A(\fifo0.fifo_data[5] ),
    .B(_03819_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_4 _07511_ (.A(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__buf_4 _07512_ (.A(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__a22o_1 _07513_ (.A1(\fifo0.fifo_store[0][5] ),
    .A2(_03827_),
    .B1(_03839_),
    .B2(_03830_),
    .X(_00012_));
 sky130_fd_sc_hd__and2_1 _07514_ (.A(\fifo0.fifo_data[6] ),
    .B(_03819_),
    .X(_03840_));
 sky130_fd_sc_hd__buf_4 _07515_ (.A(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__a22o_1 _07516_ (.A1(\fifo0.fifo_store[0][6] ),
    .A2(_03827_),
    .B1(_03841_),
    .B2(_03830_),
    .X(_00013_));
 sky130_fd_sc_hd__and2_2 _07517_ (.A(\fifo0.fifo_data[7] ),
    .B(_03819_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_4 _07518_ (.A(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__buf_4 _07519_ (.A(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__a22o_1 _07520_ (.A1(\fifo0.fifo_store[0][7] ),
    .A2(_03827_),
    .B1(_03844_),
    .B2(_03830_),
    .X(_00014_));
 sky130_fd_sc_hd__and2_1 _07521_ (.A(\fifo0.fifo_data[8] ),
    .B(_03819_),
    .X(_03845_));
 sky130_fd_sc_hd__buf_4 _07522_ (.A(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__a22o_1 _07523_ (.A1(\fifo0.fifo_store[0][8] ),
    .A2(_03827_),
    .B1(_03846_),
    .B2(_03830_),
    .X(_00015_));
 sky130_fd_sc_hd__and2_1 _07524_ (.A(\fifo0.fifo_data[9] ),
    .B(_03819_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_4 _07525_ (.A(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__a22o_1 _07526_ (.A1(\fifo0.fifo_store[0][9] ),
    .A2(_03827_),
    .B1(_03848_),
    .B2(_03830_),
    .X(_00016_));
 sky130_fd_sc_hd__and2_1 _07527_ (.A(\fifo0.fifo_data[10] ),
    .B(_03818_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_4 _07528_ (.A(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_4 _07529_ (.A(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__a22o_1 _07530_ (.A1(\fifo0.fifo_store[0][10] ),
    .A2(_03826_),
    .B1(_03851_),
    .B2(_03830_),
    .X(_00017_));
 sky130_fd_sc_hd__and2_2 _07531_ (.A(\fifo0.fifo_data[11] ),
    .B(_03818_),
    .X(_03852_));
 sky130_fd_sc_hd__buf_4 _07532_ (.A(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_4 _07533_ (.A(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__a22o_1 _07534_ (.A1(\fifo0.fifo_store[0][11] ),
    .A2(_03826_),
    .B1(_03854_),
    .B2(_03817_),
    .X(_00018_));
 sky130_fd_sc_hd__and2_1 _07535_ (.A(\fifo0.fifo_data[12] ),
    .B(_03818_),
    .X(_03855_));
 sky130_fd_sc_hd__buf_4 _07536_ (.A(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__a22o_1 _07537_ (.A1(\fifo0.fifo_store[0][12] ),
    .A2(_03826_),
    .B1(_03856_),
    .B2(_03817_),
    .X(_00019_));
 sky130_fd_sc_hd__and2_1 _07538_ (.A(\fifo0.fifo_data[13] ),
    .B(_03818_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_4 _07539_ (.A(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__a22o_1 _07540_ (.A1(\fifo0.fifo_store[0][13] ),
    .A2(_03826_),
    .B1(_03858_),
    .B2(_03817_),
    .X(_00020_));
 sky130_fd_sc_hd__and2_1 _07541_ (.A(\fifo0.fifo_data[14] ),
    .B(_03818_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_4 _07542_ (.A(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__a22o_1 _07543_ (.A1(\fifo0.fifo_store[0][14] ),
    .A2(_03826_),
    .B1(_03860_),
    .B2(_03817_),
    .X(_00021_));
 sky130_fd_sc_hd__or2_2 _07544_ (.A(\fifo0.fifo_data[15] ),
    .B(_03802_),
    .X(_03861_));
 sky130_fd_sc_hd__buf_4 _07545_ (.A(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__inv_2 _07546_ (.A(_03826_),
    .Y(_03863_));
 sky130_fd_sc_hd__o32a_1 _07547_ (.A1(_03814_),
    .A2(_03816_),
    .A3(_03862_),
    .B1(_03863_),
    .B2(\fifo0.fifo_store[0][15] ),
    .X(_00022_));
 sky130_fd_sc_hd__buf_4 _07548_ (.A(_03821_),
    .X(_03864_));
 sky130_fd_sc_hd__nand2_2 _07549_ (.A(_03803_),
    .B(_03805_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand2_2 _07550_ (.A(_03808_),
    .B(_03811_),
    .Y(_03866_));
 sky130_fd_sc_hd__or2_1 _07551_ (.A(_03865_),
    .B(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__buf_12 _07552_ (.A(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__nor2_8 _07553_ (.A(_03816_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__buf_6 _07554_ (.A(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _07555_ (.A0(\fifo0.fifo_store[80][0] ),
    .A1(_03864_),
    .S(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _07556_ (.A(_03871_),
    .X(_00023_));
 sky130_fd_sc_hd__clkbuf_4 _07557_ (.A(_03828_),
    .X(_03872_));
 sky130_fd_sc_hd__clkbuf_4 _07558_ (.A(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _07559_ (.A0(\fifo0.fifo_store[80][1] ),
    .A1(_03873_),
    .S(_03870_),
    .X(_03874_));
 sky130_fd_sc_hd__clkbuf_1 _07560_ (.A(_03874_),
    .X(_00024_));
 sky130_fd_sc_hd__clkbuf_4 _07561_ (.A(_03831_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_4 _07562_ (.A(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _07563_ (.A0(\fifo0.fifo_store[80][2] ),
    .A1(_03876_),
    .S(_03870_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _07564_ (.A(_03877_),
    .X(_00025_));
 sky130_fd_sc_hd__clkbuf_4 _07565_ (.A(_03833_),
    .X(_03878_));
 sky130_fd_sc_hd__clkbuf_4 _07566_ (.A(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__mux2_1 _07567_ (.A0(\fifo0.fifo_store[80][3] ),
    .A1(_03879_),
    .S(_03870_),
    .X(_03880_));
 sky130_fd_sc_hd__clkbuf_1 _07568_ (.A(_03880_),
    .X(_00026_));
 sky130_fd_sc_hd__clkbuf_4 _07569_ (.A(_03835_),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_4 _07570_ (.A(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__mux2_1 _07571_ (.A0(\fifo0.fifo_store[80][4] ),
    .A1(_03882_),
    .S(_03870_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _07572_ (.A(_03883_),
    .X(_00027_));
 sky130_fd_sc_hd__clkbuf_8 _07573_ (.A(_03837_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_4 _07574_ (.A(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__mux2_1 _07575_ (.A0(\fifo0.fifo_store[80][5] ),
    .A1(_03885_),
    .S(_03870_),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_1 _07576_ (.A(_03886_),
    .X(_00028_));
 sky130_fd_sc_hd__clkbuf_4 _07577_ (.A(_03840_),
    .X(_03887_));
 sky130_fd_sc_hd__buf_4 _07578_ (.A(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _07579_ (.A0(\fifo0.fifo_store[80][6] ),
    .A1(_03888_),
    .S(_03870_),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_1 _07580_ (.A(_03889_),
    .X(_00029_));
 sky130_fd_sc_hd__buf_4 _07581_ (.A(_03842_),
    .X(_03890_));
 sky130_fd_sc_hd__buf_2 _07582_ (.A(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__mux2_1 _07583_ (.A0(\fifo0.fifo_store[80][7] ),
    .A1(_03891_),
    .S(_03870_),
    .X(_03892_));
 sky130_fd_sc_hd__clkbuf_1 _07584_ (.A(_03892_),
    .X(_00030_));
 sky130_fd_sc_hd__clkbuf_4 _07585_ (.A(_03845_),
    .X(_03893_));
 sky130_fd_sc_hd__buf_2 _07586_ (.A(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__mux2_1 _07587_ (.A0(\fifo0.fifo_store[80][8] ),
    .A1(_03894_),
    .S(_03870_),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_1 _07588_ (.A(_03895_),
    .X(_00031_));
 sky130_fd_sc_hd__clkbuf_4 _07589_ (.A(_03847_),
    .X(_03896_));
 sky130_fd_sc_hd__buf_4 _07590_ (.A(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__mux2_1 _07591_ (.A0(\fifo0.fifo_store[80][9] ),
    .A1(_03897_),
    .S(_03870_),
    .X(_03898_));
 sky130_fd_sc_hd__clkbuf_1 _07592_ (.A(_03898_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_4 _07593_ (.A(_03849_),
    .X(_03899_));
 sky130_fd_sc_hd__clkbuf_4 _07594_ (.A(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _07595_ (.A0(\fifo0.fifo_store[80][10] ),
    .A1(_03900_),
    .S(_03869_),
    .X(_03901_));
 sky130_fd_sc_hd__clkbuf_1 _07596_ (.A(_03901_),
    .X(_00033_));
 sky130_fd_sc_hd__buf_6 _07597_ (.A(_03852_),
    .X(_03902_));
 sky130_fd_sc_hd__clkbuf_4 _07598_ (.A(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__mux2_1 _07599_ (.A0(\fifo0.fifo_store[80][11] ),
    .A1(_03903_),
    .S(_03869_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_1 _07600_ (.A(_03904_),
    .X(_00034_));
 sky130_fd_sc_hd__clkbuf_4 _07601_ (.A(_03855_),
    .X(_03905_));
 sky130_fd_sc_hd__buf_4 _07602_ (.A(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__mux2_1 _07603_ (.A0(\fifo0.fifo_store[80][12] ),
    .A1(_03906_),
    .S(_03869_),
    .X(_03907_));
 sky130_fd_sc_hd__clkbuf_1 _07604_ (.A(_03907_),
    .X(_00035_));
 sky130_fd_sc_hd__buf_4 _07605_ (.A(_03857_),
    .X(_03908_));
 sky130_fd_sc_hd__clkbuf_4 _07606_ (.A(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _07607_ (.A0(\fifo0.fifo_store[80][13] ),
    .A1(_03909_),
    .S(_03869_),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_1 _07608_ (.A(_03910_),
    .X(_00036_));
 sky130_fd_sc_hd__clkbuf_4 _07609_ (.A(_03859_),
    .X(_03911_));
 sky130_fd_sc_hd__buf_4 _07610_ (.A(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__mux2_1 _07611_ (.A0(\fifo0.fifo_store[80][14] ),
    .A1(_03912_),
    .S(_03869_),
    .X(_03913_));
 sky130_fd_sc_hd__clkbuf_1 _07612_ (.A(_03913_),
    .X(_00037_));
 sky130_fd_sc_hd__clkbuf_4 _07613_ (.A(_03861_),
    .X(_03914_));
 sky130_fd_sc_hd__clkbuf_4 _07614_ (.A(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _07615_ (.A0(\fifo0.fifo_store[80][15] ),
    .A1(_03915_),
    .S(_03869_),
    .X(_03916_));
 sky130_fd_sc_hd__clkbuf_1 _07616_ (.A(_03916_),
    .X(_00038_));
 sky130_fd_sc_hd__or2_1 _07617_ (.A(_03787_),
    .B(_03802_),
    .X(_03917_));
 sky130_fd_sc_hd__or3_1 _07618_ (.A(\fifo0.write_ptr[0] ),
    .B(_03789_),
    .C(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__buf_12 _07619_ (.A(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__buf_12 _07620_ (.A(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__nor2_4 _07621_ (.A(_03814_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__buf_6 _07622_ (.A(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__mux2_1 _07623_ (.A0(\fifo0.fifo_store[7][0] ),
    .A1(_03864_),
    .S(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__clkbuf_1 _07624_ (.A(_03923_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(\fifo0.fifo_store[7][1] ),
    .A1(_03873_),
    .S(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__clkbuf_1 _07626_ (.A(_03924_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _07627_ (.A0(\fifo0.fifo_store[7][2] ),
    .A1(_03876_),
    .S(_03922_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_1 _07628_ (.A(_03925_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _07629_ (.A0(\fifo0.fifo_store[7][3] ),
    .A1(_03879_),
    .S(_03922_),
    .X(_03926_));
 sky130_fd_sc_hd__clkbuf_1 _07630_ (.A(_03926_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _07631_ (.A0(\fifo0.fifo_store[7][4] ),
    .A1(_03882_),
    .S(_03922_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_1 _07632_ (.A(_03927_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _07633_ (.A0(\fifo0.fifo_store[7][5] ),
    .A1(_03885_),
    .S(_03922_),
    .X(_03928_));
 sky130_fd_sc_hd__clkbuf_1 _07634_ (.A(_03928_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(\fifo0.fifo_store[7][6] ),
    .A1(_03888_),
    .S(_03922_),
    .X(_03929_));
 sky130_fd_sc_hd__clkbuf_1 _07636_ (.A(_03929_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _07637_ (.A0(\fifo0.fifo_store[7][7] ),
    .A1(_03891_),
    .S(_03922_),
    .X(_03930_));
 sky130_fd_sc_hd__clkbuf_1 _07638_ (.A(_03930_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _07639_ (.A0(\fifo0.fifo_store[7][8] ),
    .A1(_03894_),
    .S(_03922_),
    .X(_03931_));
 sky130_fd_sc_hd__clkbuf_1 _07640_ (.A(_03931_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(\fifo0.fifo_store[7][9] ),
    .A1(_03897_),
    .S(_03922_),
    .X(_03932_));
 sky130_fd_sc_hd__clkbuf_1 _07642_ (.A(_03932_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _07643_ (.A0(\fifo0.fifo_store[7][10] ),
    .A1(_03900_),
    .S(_03921_),
    .X(_03933_));
 sky130_fd_sc_hd__clkbuf_1 _07644_ (.A(_03933_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _07645_ (.A0(\fifo0.fifo_store[7][11] ),
    .A1(_03903_),
    .S(_03921_),
    .X(_03934_));
 sky130_fd_sc_hd__clkbuf_1 _07646_ (.A(_03934_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _07647_ (.A0(\fifo0.fifo_store[7][12] ),
    .A1(_03906_),
    .S(_03921_),
    .X(_03935_));
 sky130_fd_sc_hd__clkbuf_1 _07648_ (.A(_03935_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _07649_ (.A0(\fifo0.fifo_store[7][13] ),
    .A1(_03909_),
    .S(_03921_),
    .X(_03936_));
 sky130_fd_sc_hd__clkbuf_1 _07650_ (.A(_03936_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _07651_ (.A0(\fifo0.fifo_store[7][14] ),
    .A1(_03912_),
    .S(_03921_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_1 _07652_ (.A(_03937_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _07653_ (.A0(\fifo0.fifo_store[7][15] ),
    .A1(_03915_),
    .S(_03921_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_1 _07654_ (.A(_03938_),
    .X(_00054_));
 sky130_fd_sc_hd__nand2_2 _07655_ (.A(_03794_),
    .B(_03804_),
    .Y(_03939_));
 sky130_fd_sc_hd__or2_1 _07656_ (.A(_03866_),
    .B(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_16 _07657_ (.A(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__or2_1 _07658_ (.A(_03789_),
    .B(_03802_),
    .X(_03942_));
 sky130_fd_sc_hd__or4b_4 _07659_ (.A(_03785_),
    .B(_03786_),
    .C(_03942_),
    .D_N(\fifo0.write_ptr[0] ),
    .X(_03943_));
 sky130_fd_sc_hd__or2_1 _07660_ (.A(_03941_),
    .B(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_4 _07661_ (.A(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_6 _07662_ (.A(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__mux2_1 _07663_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[78][0] ),
    .S(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__clkbuf_1 _07664_ (.A(_03947_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _07665_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[78][1] ),
    .S(_03946_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_1 _07666_ (.A(_03948_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _07667_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[78][2] ),
    .S(_03946_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_1 _07668_ (.A(_03949_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _07669_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[78][3] ),
    .S(_03946_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_1 _07670_ (.A(_03950_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _07671_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[78][4] ),
    .S(_03946_),
    .X(_03951_));
 sky130_fd_sc_hd__clkbuf_1 _07672_ (.A(_03951_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[78][5] ),
    .S(_03946_),
    .X(_03952_));
 sky130_fd_sc_hd__clkbuf_1 _07674_ (.A(_03952_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _07675_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[78][6] ),
    .S(_03946_),
    .X(_03953_));
 sky130_fd_sc_hd__clkbuf_1 _07676_ (.A(_03953_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _07677_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[78][7] ),
    .S(_03946_),
    .X(_03954_));
 sky130_fd_sc_hd__clkbuf_1 _07678_ (.A(_03954_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _07679_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[78][8] ),
    .S(_03946_),
    .X(_03955_));
 sky130_fd_sc_hd__clkbuf_1 _07680_ (.A(_03955_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _07681_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[78][9] ),
    .S(_03946_),
    .X(_03956_));
 sky130_fd_sc_hd__clkbuf_1 _07682_ (.A(_03956_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _07683_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[78][10] ),
    .S(_03945_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_1 _07684_ (.A(_03957_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _07685_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[78][11] ),
    .S(_03945_),
    .X(_03958_));
 sky130_fd_sc_hd__clkbuf_1 _07686_ (.A(_03958_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _07687_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[78][12] ),
    .S(_03945_),
    .X(_03959_));
 sky130_fd_sc_hd__clkbuf_1 _07688_ (.A(_03959_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _07689_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[78][13] ),
    .S(_03945_),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_1 _07690_ (.A(_03960_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _07691_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[78][14] ),
    .S(_03945_),
    .X(_03961_));
 sky130_fd_sc_hd__clkbuf_1 _07692_ (.A(_03961_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _07693_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[78][15] ),
    .S(_03945_),
    .X(_03962_));
 sky130_fd_sc_hd__clkbuf_1 _07694_ (.A(_03962_),
    .X(_00070_));
 sky130_fd_sc_hd__or4_1 _07695_ (.A(\fifo0.write_ptr[1] ),
    .B(\fifo0.write_ptr[0] ),
    .C(_03800_),
    .D(_03942_),
    .X(_03963_));
 sky130_fd_sc_hd__buf_12 _07696_ (.A(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__buf_12 _07697_ (.A(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__nor2_8 _07698_ (.A(_03941_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__buf_8 _07699_ (.A(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _07700_ (.A0(\fifo0.fifo_store[77][0] ),
    .A1(_03864_),
    .S(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _07701_ (.A(_03968_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _07702_ (.A0(\fifo0.fifo_store[77][1] ),
    .A1(_03873_),
    .S(_03967_),
    .X(_03969_));
 sky130_fd_sc_hd__clkbuf_1 _07703_ (.A(_03969_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _07704_ (.A0(\fifo0.fifo_store[77][2] ),
    .A1(_03876_),
    .S(_03967_),
    .X(_03970_));
 sky130_fd_sc_hd__clkbuf_1 _07705_ (.A(_03970_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _07706_ (.A0(\fifo0.fifo_store[77][3] ),
    .A1(_03879_),
    .S(_03967_),
    .X(_03971_));
 sky130_fd_sc_hd__clkbuf_1 _07707_ (.A(_03971_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _07708_ (.A0(\fifo0.fifo_store[77][4] ),
    .A1(_03882_),
    .S(_03967_),
    .X(_03972_));
 sky130_fd_sc_hd__clkbuf_1 _07709_ (.A(_03972_),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _07710_ (.A0(\fifo0.fifo_store[77][5] ),
    .A1(_03885_),
    .S(_03967_),
    .X(_03973_));
 sky130_fd_sc_hd__clkbuf_1 _07711_ (.A(_03973_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _07712_ (.A0(\fifo0.fifo_store[77][6] ),
    .A1(_03888_),
    .S(_03967_),
    .X(_03974_));
 sky130_fd_sc_hd__clkbuf_1 _07713_ (.A(_03974_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _07714_ (.A0(\fifo0.fifo_store[77][7] ),
    .A1(_03891_),
    .S(_03967_),
    .X(_03975_));
 sky130_fd_sc_hd__clkbuf_1 _07715_ (.A(_03975_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _07716_ (.A0(\fifo0.fifo_store[77][8] ),
    .A1(_03894_),
    .S(_03967_),
    .X(_03976_));
 sky130_fd_sc_hd__clkbuf_1 _07717_ (.A(_03976_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _07718_ (.A0(\fifo0.fifo_store[77][9] ),
    .A1(_03897_),
    .S(_03967_),
    .X(_03977_));
 sky130_fd_sc_hd__clkbuf_1 _07719_ (.A(_03977_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _07720_ (.A0(\fifo0.fifo_store[77][10] ),
    .A1(_03900_),
    .S(_03966_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _07721_ (.A(_03978_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _07722_ (.A0(\fifo0.fifo_store[77][11] ),
    .A1(_03903_),
    .S(_03966_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _07723_ (.A(_03979_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _07724_ (.A0(\fifo0.fifo_store[77][12] ),
    .A1(_03906_),
    .S(_03966_),
    .X(_03980_));
 sky130_fd_sc_hd__clkbuf_1 _07725_ (.A(_03980_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _07726_ (.A0(\fifo0.fifo_store[77][13] ),
    .A1(_03909_),
    .S(_03966_),
    .X(_03981_));
 sky130_fd_sc_hd__clkbuf_1 _07727_ (.A(_03981_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _07728_ (.A0(\fifo0.fifo_store[77][14] ),
    .A1(_03912_),
    .S(_03966_),
    .X(_03982_));
 sky130_fd_sc_hd__clkbuf_1 _07729_ (.A(_03982_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _07730_ (.A0(\fifo0.fifo_store[77][15] ),
    .A1(_03915_),
    .S(_03966_),
    .X(_03983_));
 sky130_fd_sc_hd__clkbuf_1 _07731_ (.A(_03983_),
    .X(_00086_));
 sky130_fd_sc_hd__or4_4 _07732_ (.A(_03799_),
    .B(_03810_),
    .C(_03800_),
    .D(_03808_),
    .X(_03984_));
 sky130_fd_sc_hd__or2_1 _07733_ (.A(_03806_),
    .B(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__buf_12 _07734_ (.A(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _07735_ (.A(\fifo0.write_ptr[0] ),
    .B(_03800_),
    .Y(_03987_));
 sky130_fd_sc_hd__or3_1 _07736_ (.A(\fifo0.write_ptr[2] ),
    .B(_03917_),
    .C(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__buf_12 _07737_ (.A(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__buf_12 _07738_ (.A(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__nor2_8 _07739_ (.A(_03986_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__buf_6 _07740_ (.A(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__mux2_1 _07741_ (.A0(\fifo0.fifo_store[98][0] ),
    .A1(_03864_),
    .S(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__clkbuf_1 _07742_ (.A(_03993_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _07743_ (.A0(\fifo0.fifo_store[98][1] ),
    .A1(_03873_),
    .S(_03992_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _07744_ (.A(_03994_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _07745_ (.A0(\fifo0.fifo_store[98][2] ),
    .A1(_03876_),
    .S(_03992_),
    .X(_03995_));
 sky130_fd_sc_hd__clkbuf_1 _07746_ (.A(_03995_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _07747_ (.A0(\fifo0.fifo_store[98][3] ),
    .A1(_03879_),
    .S(_03992_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_1 _07748_ (.A(_03996_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _07749_ (.A0(\fifo0.fifo_store[98][4] ),
    .A1(_03882_),
    .S(_03992_),
    .X(_03997_));
 sky130_fd_sc_hd__clkbuf_1 _07750_ (.A(_03997_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _07751_ (.A0(\fifo0.fifo_store[98][5] ),
    .A1(_03885_),
    .S(_03992_),
    .X(_03998_));
 sky130_fd_sc_hd__clkbuf_1 _07752_ (.A(_03998_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _07753_ (.A0(\fifo0.fifo_store[98][6] ),
    .A1(_03888_),
    .S(_03992_),
    .X(_03999_));
 sky130_fd_sc_hd__clkbuf_1 _07754_ (.A(_03999_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _07755_ (.A0(\fifo0.fifo_store[98][7] ),
    .A1(_03891_),
    .S(_03992_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _07756_ (.A(_04000_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _07757_ (.A0(\fifo0.fifo_store[98][8] ),
    .A1(_03894_),
    .S(_03992_),
    .X(_04001_));
 sky130_fd_sc_hd__clkbuf_1 _07758_ (.A(_04001_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _07759_ (.A0(\fifo0.fifo_store[98][9] ),
    .A1(_03897_),
    .S(_03992_),
    .X(_04002_));
 sky130_fd_sc_hd__clkbuf_1 _07760_ (.A(_04002_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _07761_ (.A0(\fifo0.fifo_store[98][10] ),
    .A1(_03900_),
    .S(_03991_),
    .X(_04003_));
 sky130_fd_sc_hd__clkbuf_1 _07762_ (.A(_04003_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _07763_ (.A0(\fifo0.fifo_store[98][11] ),
    .A1(_03903_),
    .S(_03991_),
    .X(_04004_));
 sky130_fd_sc_hd__clkbuf_1 _07764_ (.A(_04004_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(\fifo0.fifo_store[98][12] ),
    .A1(_03906_),
    .S(_03991_),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _07766_ (.A(_04005_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _07767_ (.A0(\fifo0.fifo_store[98][13] ),
    .A1(_03909_),
    .S(_03991_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_1 _07768_ (.A(_04006_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _07769_ (.A0(\fifo0.fifo_store[98][14] ),
    .A1(_03912_),
    .S(_03991_),
    .X(_04007_));
 sky130_fd_sc_hd__clkbuf_1 _07770_ (.A(_04007_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _07771_ (.A0(\fifo0.fifo_store[98][15] ),
    .A1(_03915_),
    .S(_03991_),
    .X(_04008_));
 sky130_fd_sc_hd__clkbuf_1 _07772_ (.A(_04008_),
    .X(_00102_));
 sky130_fd_sc_hd__or3b_1 _07773_ (.A(_03942_),
    .B(_03987_),
    .C_N(_03787_),
    .X(_04009_));
 sky130_fd_sc_hd__buf_8 _07774_ (.A(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__or2_1 _07775_ (.A(_03941_),
    .B(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__buf_4 _07776_ (.A(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__buf_6 _07777_ (.A(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_1 _07778_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[76][0] ),
    .S(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _07779_ (.A(_04014_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _07780_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[76][1] ),
    .S(_04013_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_1 _07781_ (.A(_04015_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _07782_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[76][2] ),
    .S(_04013_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_1 _07783_ (.A(_04016_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _07784_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[76][3] ),
    .S(_04013_),
    .X(_04017_));
 sky130_fd_sc_hd__clkbuf_1 _07785_ (.A(_04017_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _07786_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[76][4] ),
    .S(_04013_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _07787_ (.A(_04018_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _07788_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[76][5] ),
    .S(_04013_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_1 _07789_ (.A(_04019_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _07790_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[76][6] ),
    .S(_04013_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_1 _07791_ (.A(_04020_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _07792_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[76][7] ),
    .S(_04013_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_1 _07793_ (.A(_04021_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _07794_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[76][8] ),
    .S(_04013_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _07795_ (.A(_04022_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _07796_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[76][9] ),
    .S(_04013_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_1 _07797_ (.A(_04023_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _07798_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[76][10] ),
    .S(_04012_),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_1 _07799_ (.A(_04024_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _07800_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[76][11] ),
    .S(_04012_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _07801_ (.A(_04025_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _07802_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[76][12] ),
    .S(_04012_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _07803_ (.A(_04026_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _07804_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[76][13] ),
    .S(_04012_),
    .X(_04027_));
 sky130_fd_sc_hd__clkbuf_1 _07805_ (.A(_04027_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _07806_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[76][14] ),
    .S(_04012_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _07807_ (.A(_04028_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _07808_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[76][15] ),
    .S(_04012_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_1 _07809_ (.A(_04029_),
    .X(_00118_));
 sky130_fd_sc_hd__or3b_1 _07810_ (.A(_03802_),
    .B(\fifo0.write_ptr[2] ),
    .C_N(_03786_),
    .X(_04030_));
 sky130_fd_sc_hd__buf_12 _07811_ (.A(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__buf_12 _07812_ (.A(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_8 _07813_ (.A(_03986_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__buf_6 _07814_ (.A(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__mux2_1 _07815_ (.A0(\fifo0.fifo_store[97][0] ),
    .A1(_03864_),
    .S(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _07816_ (.A(_04035_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _07817_ (.A0(\fifo0.fifo_store[97][1] ),
    .A1(_03873_),
    .S(_04034_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _07818_ (.A(_04036_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _07819_ (.A0(\fifo0.fifo_store[97][2] ),
    .A1(_03876_),
    .S(_04034_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _07820_ (.A(_04037_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _07821_ (.A0(\fifo0.fifo_store[97][3] ),
    .A1(_03879_),
    .S(_04034_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _07822_ (.A(_04038_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _07823_ (.A0(\fifo0.fifo_store[97][4] ),
    .A1(_03882_),
    .S(_04034_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_1 _07824_ (.A(_04039_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _07825_ (.A0(\fifo0.fifo_store[97][5] ),
    .A1(_03885_),
    .S(_04034_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _07826_ (.A(_04040_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _07827_ (.A0(\fifo0.fifo_store[97][6] ),
    .A1(_03888_),
    .S(_04034_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _07828_ (.A(_04041_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _07829_ (.A0(\fifo0.fifo_store[97][7] ),
    .A1(_03891_),
    .S(_04034_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _07830_ (.A(_04042_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _07831_ (.A0(\fifo0.fifo_store[97][8] ),
    .A1(_03894_),
    .S(_04034_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _07832_ (.A(_04043_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _07833_ (.A0(\fifo0.fifo_store[97][9] ),
    .A1(_03897_),
    .S(_04034_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_1 _07834_ (.A(_04044_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _07835_ (.A0(\fifo0.fifo_store[97][10] ),
    .A1(_03900_),
    .S(_04033_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _07836_ (.A(_04045_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _07837_ (.A0(\fifo0.fifo_store[97][11] ),
    .A1(_03903_),
    .S(_04033_),
    .X(_04046_));
 sky130_fd_sc_hd__clkbuf_1 _07838_ (.A(_04046_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _07839_ (.A0(\fifo0.fifo_store[97][12] ),
    .A1(_03906_),
    .S(_04033_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _07840_ (.A(_04047_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _07841_ (.A0(\fifo0.fifo_store[97][13] ),
    .A1(_03909_),
    .S(_04033_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _07842_ (.A(_04048_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _07843_ (.A0(\fifo0.fifo_store[97][14] ),
    .A1(_03912_),
    .S(_04033_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _07844_ (.A(_04049_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _07845_ (.A0(\fifo0.fifo_store[97][15] ),
    .A1(_03915_),
    .S(_04033_),
    .X(_04050_));
 sky130_fd_sc_hd__clkbuf_1 _07846_ (.A(_04050_),
    .X(_00134_));
 sky130_fd_sc_hd__or3b_1 _07847_ (.A(\fifo0.write_ptr[2] ),
    .B(_03917_),
    .C_N(_03987_),
    .X(_04051_));
 sky130_fd_sc_hd__buf_12 _07848_ (.A(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__buf_12 _07849_ (.A(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_8 _07850_ (.A(_03941_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__clkbuf_16 _07851_ (.A(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _07852_ (.A0(\fifo0.fifo_store[75][0] ),
    .A1(_03864_),
    .S(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _07853_ (.A(_04056_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _07854_ (.A0(\fifo0.fifo_store[75][1] ),
    .A1(_03873_),
    .S(_04055_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _07855_ (.A(_04057_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _07856_ (.A0(\fifo0.fifo_store[75][2] ),
    .A1(_03876_),
    .S(_04055_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _07857_ (.A(_04058_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _07858_ (.A0(\fifo0.fifo_store[75][3] ),
    .A1(_03879_),
    .S(_04055_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_1 _07859_ (.A(_04059_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _07860_ (.A0(\fifo0.fifo_store[75][4] ),
    .A1(_03882_),
    .S(_04055_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _07861_ (.A(_04060_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _07862_ (.A0(\fifo0.fifo_store[75][5] ),
    .A1(_03885_),
    .S(_04055_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_1 _07863_ (.A(_04061_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _07864_ (.A0(\fifo0.fifo_store[75][6] ),
    .A1(_03888_),
    .S(_04055_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _07865_ (.A(_04062_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _07866_ (.A0(\fifo0.fifo_store[75][7] ),
    .A1(_03891_),
    .S(_04055_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _07867_ (.A(_04063_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _07868_ (.A0(\fifo0.fifo_store[75][8] ),
    .A1(_03894_),
    .S(_04055_),
    .X(_04064_));
 sky130_fd_sc_hd__clkbuf_1 _07869_ (.A(_04064_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _07870_ (.A0(\fifo0.fifo_store[75][9] ),
    .A1(_03897_),
    .S(_04055_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _07871_ (.A(_04065_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _07872_ (.A0(\fifo0.fifo_store[75][10] ),
    .A1(_03900_),
    .S(_04054_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _07873_ (.A(_04066_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _07874_ (.A0(\fifo0.fifo_store[75][11] ),
    .A1(_03903_),
    .S(_04054_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _07875_ (.A(_04067_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _07876_ (.A0(\fifo0.fifo_store[75][12] ),
    .A1(_03906_),
    .S(_04054_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _07877_ (.A(_04068_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _07878_ (.A0(\fifo0.fifo_store[75][13] ),
    .A1(_03909_),
    .S(_04054_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _07879_ (.A(_04069_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(\fifo0.fifo_store[75][14] ),
    .A1(_03912_),
    .S(_04054_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _07881_ (.A(_04070_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _07882_ (.A0(\fifo0.fifo_store[75][15] ),
    .A1(_03915_),
    .S(_04054_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _07883_ (.A(_04071_),
    .X(_00150_));
 sky130_fd_sc_hd__nor2_8 _07884_ (.A(_03816_),
    .B(_03986_),
    .Y(_04072_));
 sky130_fd_sc_hd__buf_6 _07885_ (.A(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__mux2_1 _07886_ (.A0(\fifo0.fifo_store[96][0] ),
    .A1(_03864_),
    .S(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _07887_ (.A(_04074_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _07888_ (.A0(\fifo0.fifo_store[96][1] ),
    .A1(_03873_),
    .S(_04073_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _07889_ (.A(_04075_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _07890_ (.A0(\fifo0.fifo_store[96][2] ),
    .A1(_03876_),
    .S(_04073_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _07891_ (.A(_04076_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _07892_ (.A0(\fifo0.fifo_store[96][3] ),
    .A1(_03879_),
    .S(_04073_),
    .X(_04077_));
 sky130_fd_sc_hd__clkbuf_1 _07893_ (.A(_04077_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _07894_ (.A0(\fifo0.fifo_store[96][4] ),
    .A1(_03882_),
    .S(_04073_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _07895_ (.A(_04078_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _07896_ (.A0(\fifo0.fifo_store[96][5] ),
    .A1(_03885_),
    .S(_04073_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _07897_ (.A(_04079_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _07898_ (.A0(\fifo0.fifo_store[96][6] ),
    .A1(_03888_),
    .S(_04073_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _07899_ (.A(_04080_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _07900_ (.A0(\fifo0.fifo_store[96][7] ),
    .A1(_03891_),
    .S(_04073_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _07901_ (.A(_04081_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _07902_ (.A0(\fifo0.fifo_store[96][8] ),
    .A1(_03894_),
    .S(_04073_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _07903_ (.A(_04082_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _07904_ (.A0(\fifo0.fifo_store[96][9] ),
    .A1(_03897_),
    .S(_04073_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _07905_ (.A(_04083_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _07906_ (.A0(\fifo0.fifo_store[96][10] ),
    .A1(_03900_),
    .S(_04072_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _07907_ (.A(_04084_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _07908_ (.A0(\fifo0.fifo_store[96][11] ),
    .A1(_03903_),
    .S(_04072_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _07909_ (.A(_04085_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _07910_ (.A0(\fifo0.fifo_store[96][12] ),
    .A1(_03906_),
    .S(_04072_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _07911_ (.A(_04086_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _07912_ (.A0(\fifo0.fifo_store[96][13] ),
    .A1(_03909_),
    .S(_04072_),
    .X(_04087_));
 sky130_fd_sc_hd__clkbuf_1 _07913_ (.A(_04087_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _07914_ (.A0(\fifo0.fifo_store[96][14] ),
    .A1(_03912_),
    .S(_04072_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _07915_ (.A(_04088_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _07916_ (.A0(\fifo0.fifo_store[96][15] ),
    .A1(_03915_),
    .S(_04072_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _07917_ (.A(_04089_),
    .X(_00166_));
 sky130_fd_sc_hd__nor2_8 _07918_ (.A(_03941_),
    .B(_03990_),
    .Y(_04090_));
 sky130_fd_sc_hd__buf_8 _07919_ (.A(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _07920_ (.A0(\fifo0.fifo_store[74][0] ),
    .A1(_03864_),
    .S(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _07921_ (.A(_04092_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _07922_ (.A0(\fifo0.fifo_store[74][1] ),
    .A1(_03873_),
    .S(_04091_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _07923_ (.A(_04093_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _07924_ (.A0(\fifo0.fifo_store[74][2] ),
    .A1(_03876_),
    .S(_04091_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _07925_ (.A(_04094_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _07926_ (.A0(\fifo0.fifo_store[74][3] ),
    .A1(_03879_),
    .S(_04091_),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _07927_ (.A(_04095_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _07928_ (.A0(\fifo0.fifo_store[74][4] ),
    .A1(_03882_),
    .S(_04091_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _07929_ (.A(_04096_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _07930_ (.A0(\fifo0.fifo_store[74][5] ),
    .A1(_03885_),
    .S(_04091_),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_1 _07931_ (.A(_04097_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _07932_ (.A0(\fifo0.fifo_store[74][6] ),
    .A1(_03888_),
    .S(_04091_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _07933_ (.A(_04098_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _07934_ (.A0(\fifo0.fifo_store[74][7] ),
    .A1(_03891_),
    .S(_04091_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _07935_ (.A(_04099_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _07936_ (.A0(\fifo0.fifo_store[74][8] ),
    .A1(_03894_),
    .S(_04091_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _07937_ (.A(_04100_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _07938_ (.A0(\fifo0.fifo_store[74][9] ),
    .A1(_03897_),
    .S(_04091_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _07939_ (.A(_04101_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _07940_ (.A0(\fifo0.fifo_store[74][10] ),
    .A1(_03900_),
    .S(_04090_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _07941_ (.A(_04102_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _07942_ (.A0(\fifo0.fifo_store[74][11] ),
    .A1(_03903_),
    .S(_04090_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _07943_ (.A(_04103_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _07944_ (.A0(\fifo0.fifo_store[74][12] ),
    .A1(_03906_),
    .S(_04090_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _07945_ (.A(_04104_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _07946_ (.A0(\fifo0.fifo_store[74][13] ),
    .A1(_03909_),
    .S(_04090_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _07947_ (.A(_04105_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _07948_ (.A0(\fifo0.fifo_store[74][14] ),
    .A1(_03912_),
    .S(_04090_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _07949_ (.A(_04106_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _07950_ (.A0(\fifo0.fifo_store[74][15] ),
    .A1(_03915_),
    .S(_04090_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _07951_ (.A(_04107_),
    .X(_00182_));
 sky130_fd_sc_hd__nor2_8 _07952_ (.A(_03941_),
    .B(_04032_),
    .Y(_04108_));
 sky130_fd_sc_hd__buf_8 _07953_ (.A(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__mux2_1 _07954_ (.A0(\fifo0.fifo_store[73][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _07955_ (.A(_04110_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _07956_ (.A0(\fifo0.fifo_store[73][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_04109_),
    .X(_04111_));
 sky130_fd_sc_hd__clkbuf_1 _07957_ (.A(_04111_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _07958_ (.A0(\fifo0.fifo_store[73][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_04109_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _07959_ (.A(_04112_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(\fifo0.fifo_store[73][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_04109_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _07961_ (.A(_04113_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _07962_ (.A0(\fifo0.fifo_store[73][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_04109_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _07963_ (.A(_04114_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _07964_ (.A0(\fifo0.fifo_store[73][5] ),
    .A1(_03885_),
    .S(_04109_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _07965_ (.A(_04115_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _07966_ (.A0(\fifo0.fifo_store[73][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_04109_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _07967_ (.A(_04116_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _07968_ (.A0(\fifo0.fifo_store[73][7] ),
    .A1(_03891_),
    .S(_04109_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _07969_ (.A(_04117_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _07970_ (.A0(\fifo0.fifo_store[73][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_04109_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _07971_ (.A(_04118_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _07972_ (.A0(\fifo0.fifo_store[73][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_04109_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _07973_ (.A(_04119_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _07974_ (.A0(\fifo0.fifo_store[73][10] ),
    .A1(_03900_),
    .S(_04108_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _07975_ (.A(_04120_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _07976_ (.A0(\fifo0.fifo_store[73][11] ),
    .A1(_03903_),
    .S(_04108_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _07977_ (.A(_04121_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _07978_ (.A0(\fifo0.fifo_store[73][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_04108_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _07979_ (.A(_04122_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _07980_ (.A0(\fifo0.fifo_store[73][13] ),
    .A1(_03909_),
    .S(_04108_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _07981_ (.A(_04123_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _07982_ (.A0(\fifo0.fifo_store[73][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_04108_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _07983_ (.A(_04124_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _07984_ (.A0(\fifo0.fifo_store[73][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_04108_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _07985_ (.A(_04125_),
    .X(_00198_));
 sky130_fd_sc_hd__nor2_8 _07986_ (.A(_03816_),
    .B(_03941_),
    .Y(_04126_));
 sky130_fd_sc_hd__buf_8 _07987_ (.A(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _07988_ (.A0(\fifo0.fifo_store[72][0] ),
    .A1(_03864_),
    .S(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _07989_ (.A(_04128_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _07990_ (.A0(\fifo0.fifo_store[72][1] ),
    .A1(_03873_),
    .S(_04127_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _07991_ (.A(_04129_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _07992_ (.A0(\fifo0.fifo_store[72][2] ),
    .A1(_03876_),
    .S(_04127_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _07993_ (.A(_04130_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _07994_ (.A0(\fifo0.fifo_store[72][3] ),
    .A1(_03879_),
    .S(_04127_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _07995_ (.A(_04131_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _07996_ (.A0(\fifo0.fifo_store[72][4] ),
    .A1(_03882_),
    .S(_04127_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _07997_ (.A(_04132_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _07998_ (.A0(\fifo0.fifo_store[72][5] ),
    .A1(_03885_),
    .S(_04127_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _07999_ (.A(_04133_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _08000_ (.A0(\fifo0.fifo_store[72][6] ),
    .A1(_03888_),
    .S(_04127_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _08001_ (.A(_04134_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _08002_ (.A0(\fifo0.fifo_store[72][7] ),
    .A1(_03891_),
    .S(_04127_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _08003_ (.A(_04135_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _08004_ (.A0(\fifo0.fifo_store[72][8] ),
    .A1(_03894_),
    .S(_04127_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _08005_ (.A(_04136_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _08006_ (.A0(\fifo0.fifo_store[72][9] ),
    .A1(_03897_),
    .S(_04127_),
    .X(_04137_));
 sky130_fd_sc_hd__clkbuf_1 _08007_ (.A(_04137_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _08008_ (.A0(\fifo0.fifo_store[72][10] ),
    .A1(_03900_),
    .S(_04126_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _08009_ (.A(_04138_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _08010_ (.A0(\fifo0.fifo_store[72][11] ),
    .A1(_03903_),
    .S(_04126_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _08011_ (.A(_04139_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _08012_ (.A0(\fifo0.fifo_store[72][12] ),
    .A1(_03906_),
    .S(_04126_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _08013_ (.A(_04140_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _08014_ (.A0(\fifo0.fifo_store[72][13] ),
    .A1(_03909_),
    .S(_04126_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _08015_ (.A(_04141_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _08016_ (.A0(\fifo0.fifo_store[72][14] ),
    .A1(_03912_),
    .S(_04126_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _08017_ (.A(_04142_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _08018_ (.A0(\fifo0.fifo_store[72][15] ),
    .A1(_03915_),
    .S(_04126_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _08019_ (.A(_04143_),
    .X(_00214_));
 sky130_fd_sc_hd__or2_1 _08020_ (.A(_03806_),
    .B(_03866_),
    .X(_04144_));
 sky130_fd_sc_hd__buf_8 _08021_ (.A(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__nor2_8 _08022_ (.A(_03920_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__buf_8 _08023_ (.A(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__mux2_1 _08024_ (.A0(\fifo0.fifo_store[71][0] ),
    .A1(_03864_),
    .S(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _08025_ (.A(_04148_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _08026_ (.A0(\fifo0.fifo_store[71][1] ),
    .A1(_03873_),
    .S(_04147_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _08027_ (.A(_04149_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _08028_ (.A0(\fifo0.fifo_store[71][2] ),
    .A1(_03876_),
    .S(_04147_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _08029_ (.A(_04150_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _08030_ (.A0(\fifo0.fifo_store[71][3] ),
    .A1(_03879_),
    .S(_04147_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _08031_ (.A(_04151_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _08032_ (.A0(\fifo0.fifo_store[71][4] ),
    .A1(_03882_),
    .S(_04147_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _08033_ (.A(_04152_),
    .X(_00219_));
 sky130_fd_sc_hd__clkbuf_4 _08034_ (.A(_03884_),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_1 _08035_ (.A0(\fifo0.fifo_store[71][5] ),
    .A1(_04153_),
    .S(_04147_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _08036_ (.A(_04154_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _08037_ (.A0(\fifo0.fifo_store[71][6] ),
    .A1(_03888_),
    .S(_04147_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _08038_ (.A(_04155_),
    .X(_00221_));
 sky130_fd_sc_hd__clkbuf_4 _08039_ (.A(_03890_),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _08040_ (.A0(\fifo0.fifo_store[71][7] ),
    .A1(_04156_),
    .S(_04147_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _08041_ (.A(_04157_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _08042_ (.A0(\fifo0.fifo_store[71][8] ),
    .A1(_03894_),
    .S(_04147_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _08043_ (.A(_04158_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _08044_ (.A0(\fifo0.fifo_store[71][9] ),
    .A1(_03897_),
    .S(_04147_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _08045_ (.A(_04159_),
    .X(_00224_));
 sky130_fd_sc_hd__clkbuf_4 _08046_ (.A(_03899_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _08047_ (.A0(\fifo0.fifo_store[71][10] ),
    .A1(_04160_),
    .S(_04146_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _08048_ (.A(_04161_),
    .X(_00225_));
 sky130_fd_sc_hd__buf_4 _08049_ (.A(_03902_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _08050_ (.A0(\fifo0.fifo_store[71][11] ),
    .A1(_04162_),
    .S(_04146_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _08051_ (.A(_04163_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _08052_ (.A0(\fifo0.fifo_store[71][12] ),
    .A1(_03906_),
    .S(_04146_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _08053_ (.A(_04164_),
    .X(_00227_));
 sky130_fd_sc_hd__buf_4 _08054_ (.A(_03908_),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _08055_ (.A0(\fifo0.fifo_store[71][13] ),
    .A1(_04165_),
    .S(_04146_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _08056_ (.A(_04166_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _08057_ (.A0(\fifo0.fifo_store[71][14] ),
    .A1(_03912_),
    .S(_04146_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _08058_ (.A(_04167_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _08059_ (.A0(\fifo0.fifo_store[71][15] ),
    .A1(_03915_),
    .S(_04146_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _08060_ (.A(_04168_),
    .X(_00230_));
 sky130_fd_sc_hd__clkbuf_4 _08061_ (.A(_03821_),
    .X(_04169_));
 sky130_fd_sc_hd__or3_2 _08062_ (.A(_03794_),
    .B(_03802_),
    .C(_03803_),
    .X(_04170_));
 sky130_fd_sc_hd__or2_2 _08063_ (.A(_03866_),
    .B(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__buf_12 _08064_ (.A(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__nor2_8 _08065_ (.A(_03920_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__buf_8 _08066_ (.A(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(\fifo0.fifo_store[95][0] ),
    .A1(_04169_),
    .S(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _08068_ (.A(_04175_),
    .X(_00231_));
 sky130_fd_sc_hd__buf_2 _08069_ (.A(_03872_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _08070_ (.A0(\fifo0.fifo_store[95][1] ),
    .A1(_04176_),
    .S(_04174_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _08071_ (.A(_04177_),
    .X(_00232_));
 sky130_fd_sc_hd__clkbuf_4 _08072_ (.A(_03875_),
    .X(_04178_));
 sky130_fd_sc_hd__mux2_1 _08073_ (.A0(\fifo0.fifo_store[95][2] ),
    .A1(_04178_),
    .S(_04174_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _08074_ (.A(_04179_),
    .X(_00233_));
 sky130_fd_sc_hd__buf_2 _08075_ (.A(_03878_),
    .X(_04180_));
 sky130_fd_sc_hd__mux2_1 _08076_ (.A0(\fifo0.fifo_store[95][3] ),
    .A1(_04180_),
    .S(_04174_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _08077_ (.A(_04181_),
    .X(_00234_));
 sky130_fd_sc_hd__buf_2 _08078_ (.A(_03881_),
    .X(_04182_));
 sky130_fd_sc_hd__mux2_1 _08079_ (.A0(\fifo0.fifo_store[95][4] ),
    .A1(_04182_),
    .S(_04174_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _08080_ (.A(_04183_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _08081_ (.A0(\fifo0.fifo_store[95][5] ),
    .A1(_04153_),
    .S(_04174_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _08082_ (.A(_04184_),
    .X(_00236_));
 sky130_fd_sc_hd__clkbuf_4 _08083_ (.A(_03887_),
    .X(_04185_));
 sky130_fd_sc_hd__mux2_1 _08084_ (.A0(\fifo0.fifo_store[95][6] ),
    .A1(_04185_),
    .S(_04174_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _08085_ (.A(_04186_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _08086_ (.A0(\fifo0.fifo_store[95][7] ),
    .A1(_04156_),
    .S(_04174_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _08087_ (.A(_04187_),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_4 _08088_ (.A(_03893_),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _08089_ (.A0(\fifo0.fifo_store[95][8] ),
    .A1(_04188_),
    .S(_04174_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _08090_ (.A(_04189_),
    .X(_00239_));
 sky130_fd_sc_hd__clkbuf_4 _08091_ (.A(_03896_),
    .X(_04190_));
 sky130_fd_sc_hd__mux2_1 _08092_ (.A0(\fifo0.fifo_store[95][9] ),
    .A1(_04190_),
    .S(_04174_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _08093_ (.A(_04191_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _08094_ (.A0(\fifo0.fifo_store[95][10] ),
    .A1(_04160_),
    .S(_04173_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _08095_ (.A(_04192_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _08096_ (.A0(\fifo0.fifo_store[95][11] ),
    .A1(_04162_),
    .S(_04173_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _08097_ (.A(_04193_),
    .X(_00242_));
 sky130_fd_sc_hd__buf_4 _08098_ (.A(_03905_),
    .X(_04194_));
 sky130_fd_sc_hd__mux2_1 _08099_ (.A0(\fifo0.fifo_store[95][12] ),
    .A1(_04194_),
    .S(_04173_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _08100_ (.A(_04195_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _08101_ (.A0(\fifo0.fifo_store[95][13] ),
    .A1(_04165_),
    .S(_04173_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _08102_ (.A(_04196_),
    .X(_00244_));
 sky130_fd_sc_hd__buf_4 _08103_ (.A(_03911_),
    .X(_04197_));
 sky130_fd_sc_hd__mux2_1 _08104_ (.A0(\fifo0.fifo_store[95][14] ),
    .A1(_04197_),
    .S(_04173_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _08105_ (.A(_04198_),
    .X(_00245_));
 sky130_fd_sc_hd__clkbuf_4 _08106_ (.A(_03914_),
    .X(_04199_));
 sky130_fd_sc_hd__mux2_1 _08107_ (.A0(\fifo0.fifo_store[95][15] ),
    .A1(_04199_),
    .S(_04173_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _08108_ (.A(_04200_),
    .X(_00246_));
 sky130_fd_sc_hd__clkbuf_4 _08109_ (.A(_03943_),
    .X(_04201_));
 sky130_fd_sc_hd__or2_1 _08110_ (.A(_04201_),
    .B(_04145_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_4 _08111_ (.A(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__buf_8 _08112_ (.A(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _08113_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[70][0] ),
    .S(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _08114_ (.A(_04205_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _08115_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[70][1] ),
    .S(_04204_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _08116_ (.A(_04206_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _08117_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[70][2] ),
    .S(_04204_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _08118_ (.A(_04207_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _08119_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[70][3] ),
    .S(_04204_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _08120_ (.A(_04208_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _08121_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[70][4] ),
    .S(_04204_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _08122_ (.A(_04209_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _08123_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[70][5] ),
    .S(_04204_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _08124_ (.A(_04210_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[70][6] ),
    .S(_04204_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _08126_ (.A(_04211_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _08127_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[70][7] ),
    .S(_04204_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _08128_ (.A(_04212_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _08129_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[70][8] ),
    .S(_04204_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _08130_ (.A(_04213_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[70][9] ),
    .S(_04204_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _08132_ (.A(_04214_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _08133_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[70][10] ),
    .S(_04203_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _08134_ (.A(_04215_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _08135_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[70][11] ),
    .S(_04203_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _08136_ (.A(_04216_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _08137_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[70][12] ),
    .S(_04203_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _08138_ (.A(_04217_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _08139_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[70][13] ),
    .S(_04203_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _08140_ (.A(_04218_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _08141_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[70][14] ),
    .S(_04203_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _08142_ (.A(_04219_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _08143_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[70][15] ),
    .S(_04203_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _08144_ (.A(_04220_),
    .X(_00262_));
 sky130_fd_sc_hd__or2_1 _08145_ (.A(_03814_),
    .B(_03943_),
    .X(_04221_));
 sky130_fd_sc_hd__buf_4 _08146_ (.A(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__buf_6 _08147_ (.A(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__mux2_1 _08148_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[6][0] ),
    .S(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _08149_ (.A(_04224_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _08150_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[6][1] ),
    .S(_04223_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _08151_ (.A(_04225_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _08152_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[6][2] ),
    .S(_04223_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _08153_ (.A(_04226_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _08154_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[6][3] ),
    .S(_04223_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _08155_ (.A(_04227_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _08156_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[6][4] ),
    .S(_04223_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _08157_ (.A(_04228_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _08158_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[6][5] ),
    .S(_04223_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _08159_ (.A(_04229_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _08160_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[6][6] ),
    .S(_04223_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _08161_ (.A(_04230_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _08162_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[6][7] ),
    .S(_04223_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _08163_ (.A(_04231_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _08164_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[6][8] ),
    .S(_04223_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _08165_ (.A(_04232_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _08166_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[6][9] ),
    .S(_04223_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _08167_ (.A(_04233_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _08168_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[6][10] ),
    .S(_04222_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _08169_ (.A(_04234_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _08170_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[6][11] ),
    .S(_04222_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _08171_ (.A(_04235_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _08172_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[6][12] ),
    .S(_04222_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _08173_ (.A(_04236_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[6][13] ),
    .S(_04222_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _08175_ (.A(_04237_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _08176_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[6][14] ),
    .S(_04222_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _08177_ (.A(_04238_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[6][15] ),
    .S(_04222_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _08179_ (.A(_04239_),
    .X(_00278_));
 sky130_fd_sc_hd__nor2_8 _08180_ (.A(_03965_),
    .B(_04172_),
    .Y(_04240_));
 sky130_fd_sc_hd__buf_8 _08181_ (.A(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__mux2_1 _08182_ (.A0(\fifo0.fifo_store[93][0] ),
    .A1(_04169_),
    .S(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _08183_ (.A(_04242_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _08184_ (.A0(\fifo0.fifo_store[93][1] ),
    .A1(_04176_),
    .S(_04241_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _08185_ (.A(_04243_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _08186_ (.A0(\fifo0.fifo_store[93][2] ),
    .A1(_04178_),
    .S(_04241_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _08187_ (.A(_04244_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _08188_ (.A0(\fifo0.fifo_store[93][3] ),
    .A1(_04180_),
    .S(_04241_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _08189_ (.A(_04245_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _08190_ (.A0(\fifo0.fifo_store[93][4] ),
    .A1(_04182_),
    .S(_04241_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _08191_ (.A(_04246_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _08192_ (.A0(\fifo0.fifo_store[93][5] ),
    .A1(_04153_),
    .S(_04241_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _08193_ (.A(_04247_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _08194_ (.A0(\fifo0.fifo_store[93][6] ),
    .A1(_04185_),
    .S(_04241_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _08195_ (.A(_04248_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _08196_ (.A0(\fifo0.fifo_store[93][7] ),
    .A1(_04156_),
    .S(_04241_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _08197_ (.A(_04249_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _08198_ (.A0(\fifo0.fifo_store[93][8] ),
    .A1(_04188_),
    .S(_04241_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _08199_ (.A(_04250_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _08200_ (.A0(\fifo0.fifo_store[93][9] ),
    .A1(_04190_),
    .S(_04241_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _08201_ (.A(_04251_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(\fifo0.fifo_store[93][10] ),
    .A1(_04160_),
    .S(_04240_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _08203_ (.A(_04252_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _08204_ (.A0(\fifo0.fifo_store[93][11] ),
    .A1(_04162_),
    .S(_04240_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _08205_ (.A(_04253_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _08206_ (.A0(\fifo0.fifo_store[93][12] ),
    .A1(_04194_),
    .S(_04240_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _08207_ (.A(_04254_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _08208_ (.A0(\fifo0.fifo_store[93][13] ),
    .A1(_04165_),
    .S(_04240_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _08209_ (.A(_04255_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _08210_ (.A0(\fifo0.fifo_store[93][14] ),
    .A1(_04197_),
    .S(_04240_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _08211_ (.A(_04256_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _08212_ (.A0(\fifo0.fifo_store[93][15] ),
    .A1(_04199_),
    .S(_04240_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _08213_ (.A(_04257_),
    .X(_00294_));
 sky130_fd_sc_hd__or2_1 _08214_ (.A(_04010_),
    .B(_04145_),
    .X(_04258_));
 sky130_fd_sc_hd__buf_4 _08215_ (.A(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__buf_8 _08216_ (.A(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _08217_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[68][0] ),
    .S(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _08218_ (.A(_04261_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _08219_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[68][1] ),
    .S(_04260_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _08220_ (.A(_04262_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[68][2] ),
    .S(_04260_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _08222_ (.A(_04263_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _08223_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[68][3] ),
    .S(_04260_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _08224_ (.A(_04264_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _08225_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[68][4] ),
    .S(_04260_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _08226_ (.A(_04265_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _08227_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[68][5] ),
    .S(_04260_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _08228_ (.A(_04266_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _08229_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[68][6] ),
    .S(_04260_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _08230_ (.A(_04267_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _08231_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[68][7] ),
    .S(_04260_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _08232_ (.A(_04268_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _08233_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[68][8] ),
    .S(_04260_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _08234_ (.A(_04269_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _08235_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[68][9] ),
    .S(_04260_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _08236_ (.A(_04270_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _08237_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[68][10] ),
    .S(_04259_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _08238_ (.A(_04271_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[68][11] ),
    .S(_04259_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _08240_ (.A(_04272_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _08241_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[68][12] ),
    .S(_04259_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _08242_ (.A(_04273_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _08243_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[68][13] ),
    .S(_04259_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _08244_ (.A(_04274_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _08245_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[68][14] ),
    .S(_04259_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _08246_ (.A(_04275_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _08247_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[68][15] ),
    .S(_04259_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _08248_ (.A(_04276_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_12 _08249_ (.A(_04010_),
    .X(_04277_));
 sky130_fd_sc_hd__nor2_8 _08250_ (.A(_04277_),
    .B(_04172_),
    .Y(_04278_));
 sky130_fd_sc_hd__buf_8 _08251_ (.A(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__mux2_1 _08252_ (.A0(\fifo0.fifo_store[92][0] ),
    .A1(_04169_),
    .S(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _08253_ (.A(_04280_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _08254_ (.A0(\fifo0.fifo_store[92][1] ),
    .A1(_04176_),
    .S(_04279_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _08255_ (.A(_04281_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _08256_ (.A0(\fifo0.fifo_store[92][2] ),
    .A1(_04178_),
    .S(_04279_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _08257_ (.A(_04282_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(\fifo0.fifo_store[92][3] ),
    .A1(_04180_),
    .S(_04279_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _08259_ (.A(_04283_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _08260_ (.A0(\fifo0.fifo_store[92][4] ),
    .A1(_04182_),
    .S(_04279_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _08261_ (.A(_04284_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _08262_ (.A0(\fifo0.fifo_store[92][5] ),
    .A1(_04153_),
    .S(_04279_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _08263_ (.A(_04285_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _08264_ (.A0(\fifo0.fifo_store[92][6] ),
    .A1(_04185_),
    .S(_04279_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _08265_ (.A(_04286_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _08266_ (.A0(\fifo0.fifo_store[92][7] ),
    .A1(_04156_),
    .S(_04279_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _08267_ (.A(_04287_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(\fifo0.fifo_store[92][8] ),
    .A1(_04188_),
    .S(_04279_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _08269_ (.A(_04288_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _08270_ (.A0(\fifo0.fifo_store[92][9] ),
    .A1(_04190_),
    .S(_04279_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _08271_ (.A(_04289_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(\fifo0.fifo_store[92][10] ),
    .A1(_04160_),
    .S(_04278_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _08273_ (.A(_04290_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _08274_ (.A0(\fifo0.fifo_store[92][11] ),
    .A1(_04162_),
    .S(_04278_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _08275_ (.A(_04291_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(\fifo0.fifo_store[92][12] ),
    .A1(_04194_),
    .S(_04278_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _08277_ (.A(_04292_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _08278_ (.A0(\fifo0.fifo_store[92][13] ),
    .A1(_04165_),
    .S(_04278_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _08279_ (.A(_04293_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _08280_ (.A0(\fifo0.fifo_store[92][14] ),
    .A1(_04197_),
    .S(_04278_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _08281_ (.A(_04294_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _08282_ (.A0(\fifo0.fifo_store[92][15] ),
    .A1(_04199_),
    .S(_04278_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _08283_ (.A(_04295_),
    .X(_00326_));
 sky130_fd_sc_hd__or2_1 _08284_ (.A(_03939_),
    .B(_03984_),
    .X(_04296_));
 sky130_fd_sc_hd__buf_12 _08285_ (.A(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__nor2_8 _08286_ (.A(_04032_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__buf_12 _08287_ (.A(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _08288_ (.A0(\fifo0.fifo_store[105][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _08289_ (.A(_04300_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _08290_ (.A0(\fifo0.fifo_store[105][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_04299_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _08291_ (.A(_04301_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _08292_ (.A0(\fifo0.fifo_store[105][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_04299_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _08293_ (.A(_04302_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(\fifo0.fifo_store[105][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_04299_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _08295_ (.A(_04303_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _08296_ (.A0(\fifo0.fifo_store[105][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_04299_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _08297_ (.A(_04304_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(\fifo0.fifo_store[105][5] ),
    .A1(_04153_),
    .S(_04299_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _08299_ (.A(_04305_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _08300_ (.A0(\fifo0.fifo_store[105][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_04299_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _08301_ (.A(_04306_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _08302_ (.A0(\fifo0.fifo_store[105][7] ),
    .A1(_04156_),
    .S(_04299_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _08303_ (.A(_04307_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _08304_ (.A0(\fifo0.fifo_store[105][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_04299_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _08305_ (.A(_04308_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _08306_ (.A0(\fifo0.fifo_store[105][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_04299_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _08307_ (.A(_04309_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _08308_ (.A0(\fifo0.fifo_store[105][10] ),
    .A1(_04160_),
    .S(_04298_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _08309_ (.A(_04310_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _08310_ (.A0(\fifo0.fifo_store[105][11] ),
    .A1(_04162_),
    .S(_04298_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _08311_ (.A(_04311_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _08312_ (.A0(\fifo0.fifo_store[105][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_04298_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _08313_ (.A(_04312_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _08314_ (.A0(\fifo0.fifo_store[105][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_04298_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _08315_ (.A(_04313_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _08316_ (.A0(\fifo0.fifo_store[105][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_04298_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _08317_ (.A(_04314_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(\fifo0.fifo_store[105][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_04298_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _08319_ (.A(_04315_),
    .X(_00342_));
 sky130_fd_sc_hd__or2_1 _08320_ (.A(_03865_),
    .B(_03984_),
    .X(_04316_));
 sky130_fd_sc_hd__buf_8 _08321_ (.A(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__or2_1 _08322_ (.A(_04201_),
    .B(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_4 _08323_ (.A(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__buf_6 _08324_ (.A(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _08325_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[118][0] ),
    .S(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _08326_ (.A(_04321_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _08327_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[118][1] ),
    .S(_04320_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _08328_ (.A(_04322_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _08329_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[118][2] ),
    .S(_04320_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _08330_ (.A(_04323_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _08331_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[118][3] ),
    .S(_04320_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _08332_ (.A(_04324_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _08333_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[118][4] ),
    .S(_04320_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _08334_ (.A(_04325_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _08335_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[118][5] ),
    .S(_04320_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _08336_ (.A(_04326_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _08337_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[118][6] ),
    .S(_04320_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _08338_ (.A(_04327_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _08339_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[118][7] ),
    .S(_04320_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _08340_ (.A(_04328_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _08341_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[118][8] ),
    .S(_04320_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _08342_ (.A(_04329_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _08343_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[118][9] ),
    .S(_04320_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _08344_ (.A(_04330_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _08345_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[118][10] ),
    .S(_04319_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _08346_ (.A(_04331_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _08347_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[118][11] ),
    .S(_04319_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _08348_ (.A(_04332_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[118][12] ),
    .S(_04319_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _08350_ (.A(_04333_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _08351_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[118][13] ),
    .S(_04319_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _08352_ (.A(_04334_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _08353_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[118][14] ),
    .S(_04319_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _08354_ (.A(_04335_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _08355_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[118][15] ),
    .S(_04319_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _08356_ (.A(_04336_),
    .X(_00358_));
 sky130_fd_sc_hd__nor2_4 _08357_ (.A(_04053_),
    .B(_04317_),
    .Y(_04337_));
 sky130_fd_sc_hd__buf_6 _08358_ (.A(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_1 _08359_ (.A0(\fifo0.fifo_store[115][0] ),
    .A1(_04169_),
    .S(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _08360_ (.A(_04339_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _08361_ (.A0(\fifo0.fifo_store[115][1] ),
    .A1(_04176_),
    .S(_04338_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _08362_ (.A(_04340_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _08363_ (.A0(\fifo0.fifo_store[115][2] ),
    .A1(_04178_),
    .S(_04338_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _08364_ (.A(_04341_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _08365_ (.A0(\fifo0.fifo_store[115][3] ),
    .A1(_04180_),
    .S(_04338_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _08366_ (.A(_04342_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _08367_ (.A0(\fifo0.fifo_store[115][4] ),
    .A1(_04182_),
    .S(_04338_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _08368_ (.A(_04343_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _08369_ (.A0(\fifo0.fifo_store[115][5] ),
    .A1(_04153_),
    .S(_04338_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _08370_ (.A(_04344_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _08371_ (.A0(\fifo0.fifo_store[115][6] ),
    .A1(_04185_),
    .S(_04338_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _08372_ (.A(_04345_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _08373_ (.A0(\fifo0.fifo_store[115][7] ),
    .A1(_04156_),
    .S(_04338_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _08374_ (.A(_04346_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _08375_ (.A0(\fifo0.fifo_store[115][8] ),
    .A1(_04188_),
    .S(_04338_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _08376_ (.A(_04347_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _08377_ (.A0(\fifo0.fifo_store[115][9] ),
    .A1(_04190_),
    .S(_04338_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _08378_ (.A(_04348_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(\fifo0.fifo_store[115][10] ),
    .A1(_04160_),
    .S(_04337_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _08380_ (.A(_04349_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _08381_ (.A0(\fifo0.fifo_store[115][11] ),
    .A1(_04162_),
    .S(_04337_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _08382_ (.A(_04350_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _08383_ (.A0(\fifo0.fifo_store[115][12] ),
    .A1(_04194_),
    .S(_04337_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _08384_ (.A(_04351_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(\fifo0.fifo_store[115][13] ),
    .A1(_04165_),
    .S(_04337_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _08386_ (.A(_04352_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _08387_ (.A0(\fifo0.fifo_store[115][14] ),
    .A1(_04197_),
    .S(_04337_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _08388_ (.A(_04353_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(\fifo0.fifo_store[115][15] ),
    .A1(_04199_),
    .S(_04337_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _08390_ (.A(_04354_),
    .X(_00374_));
 sky130_fd_sc_hd__or2_1 _08391_ (.A(_03812_),
    .B(_03939_),
    .X(_04355_));
 sky130_fd_sc_hd__buf_12 _08392_ (.A(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__nor2_8 _08393_ (.A(_04053_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__buf_12 _08394_ (.A(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(\fifo0.fifo_store[11][0] ),
    .A1(_04169_),
    .S(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _08396_ (.A(_04359_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _08397_ (.A0(\fifo0.fifo_store[11][1] ),
    .A1(_04176_),
    .S(_04358_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _08398_ (.A(_04360_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(\fifo0.fifo_store[11][2] ),
    .A1(_04178_),
    .S(_04358_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _08400_ (.A(_04361_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _08401_ (.A0(\fifo0.fifo_store[11][3] ),
    .A1(_04180_),
    .S(_04358_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _08402_ (.A(_04362_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _08403_ (.A0(\fifo0.fifo_store[11][4] ),
    .A1(_04182_),
    .S(_04358_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _08404_ (.A(_04363_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(\fifo0.fifo_store[11][5] ),
    .A1(_04153_),
    .S(_04358_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _08406_ (.A(_04364_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _08407_ (.A0(\fifo0.fifo_store[11][6] ),
    .A1(_04185_),
    .S(_04358_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _08408_ (.A(_04365_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _08409_ (.A0(\fifo0.fifo_store[11][7] ),
    .A1(_04156_),
    .S(_04358_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _08410_ (.A(_04366_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _08411_ (.A0(\fifo0.fifo_store[11][8] ),
    .A1(_04188_),
    .S(_04358_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _08412_ (.A(_04367_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _08413_ (.A0(\fifo0.fifo_store[11][9] ),
    .A1(_04190_),
    .S(_04358_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _08414_ (.A(_04368_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(\fifo0.fifo_store[11][10] ),
    .A1(_04160_),
    .S(_04357_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _08416_ (.A(_04369_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _08417_ (.A0(\fifo0.fifo_store[11][11] ),
    .A1(_04162_),
    .S(_04357_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _08418_ (.A(_04370_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _08419_ (.A0(\fifo0.fifo_store[11][12] ),
    .A1(_04194_),
    .S(_04357_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _08420_ (.A(_04371_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _08421_ (.A0(\fifo0.fifo_store[11][13] ),
    .A1(_04165_),
    .S(_04357_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _08422_ (.A(_04372_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _08423_ (.A0(\fifo0.fifo_store[11][14] ),
    .A1(_04197_),
    .S(_04357_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _08424_ (.A(_04373_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(\fifo0.fifo_store[11][15] ),
    .A1(_04199_),
    .S(_04357_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _08426_ (.A(_04374_),
    .X(_00390_));
 sky130_fd_sc_hd__or2_1 _08427_ (.A(_03984_),
    .B(_04170_),
    .X(_04375_));
 sky130_fd_sc_hd__buf_12 _08428_ (.A(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nor2_8 _08429_ (.A(_03816_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__buf_6 _08430_ (.A(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _08431_ (.A0(\fifo0.fifo_store[120][0] ),
    .A1(_04169_),
    .S(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _08432_ (.A(_04379_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _08433_ (.A0(\fifo0.fifo_store[120][1] ),
    .A1(_04176_),
    .S(_04378_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _08434_ (.A(_04380_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(\fifo0.fifo_store[120][2] ),
    .A1(_04178_),
    .S(_04378_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _08436_ (.A(_04381_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _08437_ (.A0(\fifo0.fifo_store[120][3] ),
    .A1(_04180_),
    .S(_04378_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _08438_ (.A(_04382_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(\fifo0.fifo_store[120][4] ),
    .A1(_04182_),
    .S(_04378_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _08440_ (.A(_04383_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(\fifo0.fifo_store[120][5] ),
    .A1(_04153_),
    .S(_04378_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _08442_ (.A(_04384_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(\fifo0.fifo_store[120][6] ),
    .A1(_04185_),
    .S(_04378_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_04385_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _08445_ (.A0(\fifo0.fifo_store[120][7] ),
    .A1(_04156_),
    .S(_04378_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _08446_ (.A(_04386_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _08447_ (.A0(\fifo0.fifo_store[120][8] ),
    .A1(_04188_),
    .S(_04378_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _08448_ (.A(_04387_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _08449_ (.A0(\fifo0.fifo_store[120][9] ),
    .A1(_04190_),
    .S(_04378_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _08450_ (.A(_04388_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(\fifo0.fifo_store[120][10] ),
    .A1(_04160_),
    .S(_04377_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _08452_ (.A(_04389_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _08453_ (.A0(\fifo0.fifo_store[120][11] ),
    .A1(_04162_),
    .S(_04377_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _08454_ (.A(_04390_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _08455_ (.A0(\fifo0.fifo_store[120][12] ),
    .A1(_04194_),
    .S(_04377_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _08456_ (.A(_04391_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _08457_ (.A0(\fifo0.fifo_store[120][13] ),
    .A1(_04165_),
    .S(_04377_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _08458_ (.A(_04392_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _08459_ (.A0(\fifo0.fifo_store[120][14] ),
    .A1(_04197_),
    .S(_04377_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _08460_ (.A(_04393_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(\fifo0.fifo_store[120][15] ),
    .A1(_04199_),
    .S(_04377_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _08462_ (.A(_04394_),
    .X(_00406_));
 sky130_fd_sc_hd__nor2_8 _08463_ (.A(_04032_),
    .B(_04376_),
    .Y(_04395_));
 sky130_fd_sc_hd__buf_6 _08464_ (.A(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__mux2_1 _08465_ (.A0(\fifo0.fifo_store[121][0] ),
    .A1(_04169_),
    .S(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _08466_ (.A(_04397_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _08467_ (.A0(\fifo0.fifo_store[121][1] ),
    .A1(_04176_),
    .S(_04396_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _08468_ (.A(_04398_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _08469_ (.A0(\fifo0.fifo_store[121][2] ),
    .A1(_04178_),
    .S(_04396_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _08470_ (.A(_04399_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _08471_ (.A0(\fifo0.fifo_store[121][3] ),
    .A1(_04180_),
    .S(_04396_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _08472_ (.A(_04400_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _08473_ (.A0(\fifo0.fifo_store[121][4] ),
    .A1(_04182_),
    .S(_04396_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _08474_ (.A(_04401_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _08475_ (.A0(\fifo0.fifo_store[121][5] ),
    .A1(_04153_),
    .S(_04396_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _08476_ (.A(_04402_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _08477_ (.A0(\fifo0.fifo_store[121][6] ),
    .A1(_04185_),
    .S(_04396_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _08478_ (.A(_04403_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _08479_ (.A0(\fifo0.fifo_store[121][7] ),
    .A1(_04156_),
    .S(_04396_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _08480_ (.A(_04404_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _08481_ (.A0(\fifo0.fifo_store[121][8] ),
    .A1(_04188_),
    .S(_04396_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _08482_ (.A(_04405_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _08483_ (.A0(\fifo0.fifo_store[121][9] ),
    .A1(_04190_),
    .S(_04396_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _08484_ (.A(_04406_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _08485_ (.A0(\fifo0.fifo_store[121][10] ),
    .A1(_04160_),
    .S(_04395_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _08486_ (.A(_04407_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(\fifo0.fifo_store[121][11] ),
    .A1(_04162_),
    .S(_04395_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _08488_ (.A(_04408_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _08489_ (.A0(\fifo0.fifo_store[121][12] ),
    .A1(_04194_),
    .S(_04395_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _08490_ (.A(_04409_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(\fifo0.fifo_store[121][13] ),
    .A1(_04165_),
    .S(_04395_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _08492_ (.A(_04410_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _08493_ (.A0(\fifo0.fifo_store[121][14] ),
    .A1(_04197_),
    .S(_04395_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _08494_ (.A(_04411_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _08495_ (.A0(\fifo0.fifo_store[121][15] ),
    .A1(_04199_),
    .S(_04395_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _08496_ (.A(_04412_),
    .X(_00422_));
 sky130_fd_sc_hd__nor2_8 _08497_ (.A(_03990_),
    .B(_04376_),
    .Y(_04413_));
 sky130_fd_sc_hd__buf_6 _08498_ (.A(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__mux2_1 _08499_ (.A0(\fifo0.fifo_store[122][0] ),
    .A1(_04169_),
    .S(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _08500_ (.A(_04415_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(\fifo0.fifo_store[122][1] ),
    .A1(_04176_),
    .S(_04414_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _08502_ (.A(_04416_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(\fifo0.fifo_store[122][2] ),
    .A1(_04178_),
    .S(_04414_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _08504_ (.A(_04417_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(\fifo0.fifo_store[122][3] ),
    .A1(_04180_),
    .S(_04414_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _08506_ (.A(_04418_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(\fifo0.fifo_store[122][4] ),
    .A1(_04182_),
    .S(_04414_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _08508_ (.A(_04419_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _08509_ (.A0(\fifo0.fifo_store[122][5] ),
    .A1(_04153_),
    .S(_04414_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _08510_ (.A(_04420_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _08511_ (.A0(\fifo0.fifo_store[122][6] ),
    .A1(_04185_),
    .S(_04414_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _08512_ (.A(_04421_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _08513_ (.A0(\fifo0.fifo_store[122][7] ),
    .A1(_04156_),
    .S(_04414_),
    .X(_04422_));
 sky130_fd_sc_hd__clkbuf_1 _08514_ (.A(_04422_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _08515_ (.A0(\fifo0.fifo_store[122][8] ),
    .A1(_04188_),
    .S(_04414_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _08516_ (.A(_04423_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _08517_ (.A0(\fifo0.fifo_store[122][9] ),
    .A1(_04190_),
    .S(_04414_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _08518_ (.A(_04424_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(\fifo0.fifo_store[122][10] ),
    .A1(_04160_),
    .S(_04413_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _08520_ (.A(_04425_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _08521_ (.A0(\fifo0.fifo_store[122][11] ),
    .A1(_04162_),
    .S(_04413_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _08522_ (.A(_04426_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _08523_ (.A0(\fifo0.fifo_store[122][12] ),
    .A1(_04194_),
    .S(_04413_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _08524_ (.A(_04427_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _08525_ (.A0(\fifo0.fifo_store[122][13] ),
    .A1(_04165_),
    .S(_04413_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _08526_ (.A(_04428_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _08527_ (.A0(\fifo0.fifo_store[122][14] ),
    .A1(_04197_),
    .S(_04413_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _08528_ (.A(_04429_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _08529_ (.A0(\fifo0.fifo_store[122][15] ),
    .A1(_04199_),
    .S(_04413_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _08530_ (.A(_04430_),
    .X(_00438_));
 sky130_fd_sc_hd__nor2_4 _08531_ (.A(_04277_),
    .B(_04317_),
    .Y(_04431_));
 sky130_fd_sc_hd__buf_6 _08532_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__mux2_1 _08533_ (.A0(\fifo0.fifo_store[116][0] ),
    .A1(_04169_),
    .S(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _08534_ (.A(_04433_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(\fifo0.fifo_store[116][1] ),
    .A1(_04176_),
    .S(_04432_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _08536_ (.A(_04434_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _08537_ (.A0(\fifo0.fifo_store[116][2] ),
    .A1(_04178_),
    .S(_04432_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _08538_ (.A(_04435_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _08539_ (.A0(\fifo0.fifo_store[116][3] ),
    .A1(_04180_),
    .S(_04432_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _08540_ (.A(_04436_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _08541_ (.A0(\fifo0.fifo_store[116][4] ),
    .A1(_04182_),
    .S(_04432_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _08542_ (.A(_04437_),
    .X(_00443_));
 sky130_fd_sc_hd__clkbuf_4 _08543_ (.A(_03838_),
    .X(_04438_));
 sky130_fd_sc_hd__mux2_1 _08544_ (.A0(\fifo0.fifo_store[116][5] ),
    .A1(_04438_),
    .S(_04432_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _08545_ (.A(_04439_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(\fifo0.fifo_store[116][6] ),
    .A1(_04185_),
    .S(_04432_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _08547_ (.A(_04440_),
    .X(_00445_));
 sky130_fd_sc_hd__clkbuf_4 _08548_ (.A(_03843_),
    .X(_04441_));
 sky130_fd_sc_hd__mux2_1 _08549_ (.A0(\fifo0.fifo_store[116][7] ),
    .A1(_04441_),
    .S(_04432_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _08550_ (.A(_04442_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _08551_ (.A0(\fifo0.fifo_store[116][8] ),
    .A1(_04188_),
    .S(_04432_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _08552_ (.A(_04443_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(\fifo0.fifo_store[116][9] ),
    .A1(_04190_),
    .S(_04432_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _08554_ (.A(_04444_),
    .X(_00448_));
 sky130_fd_sc_hd__clkbuf_4 _08555_ (.A(_03850_),
    .X(_04445_));
 sky130_fd_sc_hd__mux2_1 _08556_ (.A0(\fifo0.fifo_store[116][10] ),
    .A1(_04445_),
    .S(_04431_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _08557_ (.A(_04446_),
    .X(_00449_));
 sky130_fd_sc_hd__buf_4 _08558_ (.A(_03853_),
    .X(_04447_));
 sky130_fd_sc_hd__mux2_1 _08559_ (.A0(\fifo0.fifo_store[116][11] ),
    .A1(_04447_),
    .S(_04431_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _08560_ (.A(_04448_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _08561_ (.A0(\fifo0.fifo_store[116][12] ),
    .A1(_04194_),
    .S(_04431_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _08562_ (.A(_04449_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _08563_ (.A0(\fifo0.fifo_store[116][13] ),
    .A1(_04165_),
    .S(_04431_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _08564_ (.A(_04450_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _08565_ (.A0(\fifo0.fifo_store[116][14] ),
    .A1(_04197_),
    .S(_04431_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _08566_ (.A(_04451_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _08567_ (.A0(\fifo0.fifo_store[116][15] ),
    .A1(_04199_),
    .S(_04431_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _08568_ (.A(_04452_),
    .X(_00454_));
 sky130_fd_sc_hd__nor2_8 _08569_ (.A(_04053_),
    .B(_04376_),
    .Y(_04453_));
 sky130_fd_sc_hd__buf_6 _08570_ (.A(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__mux2_1 _08571_ (.A0(\fifo0.fifo_store[123][0] ),
    .A1(_04169_),
    .S(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _08572_ (.A(_04455_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _08573_ (.A0(\fifo0.fifo_store[123][1] ),
    .A1(_04176_),
    .S(_04454_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _08574_ (.A(_04456_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _08575_ (.A0(\fifo0.fifo_store[123][2] ),
    .A1(_04178_),
    .S(_04454_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _08576_ (.A(_04457_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _08577_ (.A0(\fifo0.fifo_store[123][3] ),
    .A1(_04180_),
    .S(_04454_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _08578_ (.A(_04458_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _08579_ (.A0(\fifo0.fifo_store[123][4] ),
    .A1(_04182_),
    .S(_04454_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_1 _08580_ (.A(_04459_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _08581_ (.A0(\fifo0.fifo_store[123][5] ),
    .A1(_04438_),
    .S(_04454_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _08582_ (.A(_04460_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _08583_ (.A0(\fifo0.fifo_store[123][6] ),
    .A1(_04185_),
    .S(_04454_),
    .X(_04461_));
 sky130_fd_sc_hd__clkbuf_1 _08584_ (.A(_04461_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _08585_ (.A0(\fifo0.fifo_store[123][7] ),
    .A1(_04441_),
    .S(_04454_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _08586_ (.A(_04462_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _08587_ (.A0(\fifo0.fifo_store[123][8] ),
    .A1(_04188_),
    .S(_04454_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_1 _08588_ (.A(_04463_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _08589_ (.A0(\fifo0.fifo_store[123][9] ),
    .A1(_04190_),
    .S(_04454_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _08590_ (.A(_04464_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _08591_ (.A0(\fifo0.fifo_store[123][10] ),
    .A1(_04445_),
    .S(_04453_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _08592_ (.A(_04465_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _08593_ (.A0(\fifo0.fifo_store[123][11] ),
    .A1(_04447_),
    .S(_04453_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _08594_ (.A(_04466_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(\fifo0.fifo_store[123][12] ),
    .A1(_04194_),
    .S(_04453_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _08596_ (.A(_04467_),
    .X(_00467_));
 sky130_fd_sc_hd__buf_4 _08597_ (.A(_03908_),
    .X(_04468_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(\fifo0.fifo_store[123][13] ),
    .A1(_04468_),
    .S(_04453_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _08599_ (.A(_04469_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _08600_ (.A0(\fifo0.fifo_store[123][14] ),
    .A1(_04197_),
    .S(_04453_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _08601_ (.A(_04470_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _08602_ (.A0(\fifo0.fifo_store[123][15] ),
    .A1(_04199_),
    .S(_04453_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _08603_ (.A(_04471_),
    .X(_00470_));
 sky130_fd_sc_hd__clkbuf_4 _08604_ (.A(_03821_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_4 _08605_ (.A(_03965_),
    .B(_04317_),
    .Y(_04473_));
 sky130_fd_sc_hd__buf_6 _08606_ (.A(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _08607_ (.A0(\fifo0.fifo_store[117][0] ),
    .A1(_04472_),
    .S(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _08608_ (.A(_04475_),
    .X(_00471_));
 sky130_fd_sc_hd__clkbuf_4 _08609_ (.A(_03872_),
    .X(_04476_));
 sky130_fd_sc_hd__mux2_1 _08610_ (.A0(\fifo0.fifo_store[117][1] ),
    .A1(_04476_),
    .S(_04474_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _08611_ (.A(_04477_),
    .X(_00472_));
 sky130_fd_sc_hd__clkbuf_4 _08612_ (.A(_03875_),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(\fifo0.fifo_store[117][2] ),
    .A1(_04478_),
    .S(_04474_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _08614_ (.A(_04479_),
    .X(_00473_));
 sky130_fd_sc_hd__buf_4 _08615_ (.A(_03878_),
    .X(_04480_));
 sky130_fd_sc_hd__mux2_1 _08616_ (.A0(\fifo0.fifo_store[117][3] ),
    .A1(_04480_),
    .S(_04474_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _08617_ (.A(_04481_),
    .X(_00474_));
 sky130_fd_sc_hd__clkbuf_4 _08618_ (.A(_03881_),
    .X(_04482_));
 sky130_fd_sc_hd__mux2_1 _08619_ (.A0(\fifo0.fifo_store[117][4] ),
    .A1(_04482_),
    .S(_04474_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _08620_ (.A(_04483_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(\fifo0.fifo_store[117][5] ),
    .A1(_04438_),
    .S(_04474_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _08622_ (.A(_04484_),
    .X(_00476_));
 sky130_fd_sc_hd__clkbuf_4 _08623_ (.A(_03887_),
    .X(_04485_));
 sky130_fd_sc_hd__mux2_1 _08624_ (.A0(\fifo0.fifo_store[117][6] ),
    .A1(_04485_),
    .S(_04474_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _08625_ (.A(_04486_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _08626_ (.A0(\fifo0.fifo_store[117][7] ),
    .A1(_04441_),
    .S(_04474_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _08627_ (.A(_04487_),
    .X(_00478_));
 sky130_fd_sc_hd__buf_4 _08628_ (.A(_03893_),
    .X(_04488_));
 sky130_fd_sc_hd__mux2_1 _08629_ (.A0(\fifo0.fifo_store[117][8] ),
    .A1(_04488_),
    .S(_04474_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _08630_ (.A(_04489_),
    .X(_00479_));
 sky130_fd_sc_hd__clkbuf_4 _08631_ (.A(_03896_),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _08632_ (.A0(\fifo0.fifo_store[117][9] ),
    .A1(_04490_),
    .S(_04474_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _08633_ (.A(_04491_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _08634_ (.A0(\fifo0.fifo_store[117][10] ),
    .A1(_04445_),
    .S(_04473_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _08635_ (.A(_04492_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _08636_ (.A0(\fifo0.fifo_store[117][11] ),
    .A1(_04447_),
    .S(_04473_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _08637_ (.A(_04493_),
    .X(_00482_));
 sky130_fd_sc_hd__buf_4 _08638_ (.A(_03905_),
    .X(_04494_));
 sky130_fd_sc_hd__mux2_1 _08639_ (.A0(\fifo0.fifo_store[117][12] ),
    .A1(_04494_),
    .S(_04473_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _08640_ (.A(_04495_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _08641_ (.A0(\fifo0.fifo_store[117][13] ),
    .A1(_04468_),
    .S(_04473_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _08642_ (.A(_04496_),
    .X(_00484_));
 sky130_fd_sc_hd__buf_4 _08643_ (.A(_03911_),
    .X(_04497_));
 sky130_fd_sc_hd__mux2_1 _08644_ (.A0(\fifo0.fifo_store[117][14] ),
    .A1(_04497_),
    .S(_04473_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _08645_ (.A(_04498_),
    .X(_00485_));
 sky130_fd_sc_hd__clkbuf_4 _08646_ (.A(_03914_),
    .X(_04499_));
 sky130_fd_sc_hd__mux2_1 _08647_ (.A0(\fifo0.fifo_store[117][15] ),
    .A1(_04499_),
    .S(_04473_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _08648_ (.A(_04500_),
    .X(_00486_));
 sky130_fd_sc_hd__nor2_4 _08649_ (.A(_04277_),
    .B(_04376_),
    .Y(_04501_));
 sky130_fd_sc_hd__buf_6 _08650_ (.A(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__mux2_1 _08651_ (.A0(\fifo0.fifo_store[124][0] ),
    .A1(_04472_),
    .S(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _08652_ (.A(_04503_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _08653_ (.A0(\fifo0.fifo_store[124][1] ),
    .A1(_04476_),
    .S(_04502_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _08654_ (.A(_04504_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _08655_ (.A0(\fifo0.fifo_store[124][2] ),
    .A1(_04478_),
    .S(_04502_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_1 _08656_ (.A(_04505_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _08657_ (.A0(\fifo0.fifo_store[124][3] ),
    .A1(_04480_),
    .S(_04502_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _08658_ (.A(_04506_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _08659_ (.A0(\fifo0.fifo_store[124][4] ),
    .A1(_04482_),
    .S(_04502_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_1 _08660_ (.A(_04507_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _08661_ (.A0(\fifo0.fifo_store[124][5] ),
    .A1(_04438_),
    .S(_04502_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _08662_ (.A(_04508_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _08663_ (.A0(\fifo0.fifo_store[124][6] ),
    .A1(_04485_),
    .S(_04502_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _08664_ (.A(_04509_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _08665_ (.A0(\fifo0.fifo_store[124][7] ),
    .A1(_04441_),
    .S(_04502_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _08666_ (.A(_04510_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _08667_ (.A0(\fifo0.fifo_store[124][8] ),
    .A1(_04488_),
    .S(_04502_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _08668_ (.A(_04511_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _08669_ (.A0(\fifo0.fifo_store[124][9] ),
    .A1(_04490_),
    .S(_04502_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_1 _08670_ (.A(_04512_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _08671_ (.A0(\fifo0.fifo_store[124][10] ),
    .A1(_04445_),
    .S(_04501_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _08672_ (.A(_04513_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _08673_ (.A0(\fifo0.fifo_store[124][11] ),
    .A1(_04447_),
    .S(_04501_),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_1 _08674_ (.A(_04514_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(\fifo0.fifo_store[124][12] ),
    .A1(_04494_),
    .S(_04501_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _08676_ (.A(_04515_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(\fifo0.fifo_store[124][13] ),
    .A1(_04468_),
    .S(_04501_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _08678_ (.A(_04516_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _08679_ (.A0(\fifo0.fifo_store[124][14] ),
    .A1(_04497_),
    .S(_04501_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _08680_ (.A(_04517_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _08681_ (.A0(\fifo0.fifo_store[124][15] ),
    .A1(_04499_),
    .S(_04501_),
    .X(_04518_));
 sky130_fd_sc_hd__clkbuf_1 _08682_ (.A(_04518_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_4 _08683_ (.A(_04053_),
    .B(_04145_),
    .Y(_04519_));
 sky130_fd_sc_hd__buf_6 _08684_ (.A(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__mux2_1 _08685_ (.A0(\fifo0.fifo_store[67][0] ),
    .A1(_04472_),
    .S(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _08686_ (.A(_04521_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _08687_ (.A0(\fifo0.fifo_store[67][1] ),
    .A1(_04476_),
    .S(_04520_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _08688_ (.A(_04522_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _08689_ (.A0(\fifo0.fifo_store[67][2] ),
    .A1(_04478_),
    .S(_04520_),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_1 _08690_ (.A(_04523_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _08691_ (.A0(\fifo0.fifo_store[67][3] ),
    .A1(_04480_),
    .S(_04520_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _08692_ (.A(_04524_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _08693_ (.A0(\fifo0.fifo_store[67][4] ),
    .A1(_04482_),
    .S(_04520_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_1 _08694_ (.A(_04525_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(\fifo0.fifo_store[67][5] ),
    .A1(_04438_),
    .S(_04520_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _08696_ (.A(_04526_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _08697_ (.A0(\fifo0.fifo_store[67][6] ),
    .A1(_04485_),
    .S(_04520_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _08698_ (.A(_04527_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _08699_ (.A0(\fifo0.fifo_store[67][7] ),
    .A1(_04441_),
    .S(_04520_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _08700_ (.A(_04528_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _08701_ (.A0(\fifo0.fifo_store[67][8] ),
    .A1(_04488_),
    .S(_04520_),
    .X(_04529_));
 sky130_fd_sc_hd__clkbuf_1 _08702_ (.A(_04529_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _08703_ (.A0(\fifo0.fifo_store[67][9] ),
    .A1(_04490_),
    .S(_04520_),
    .X(_04530_));
 sky130_fd_sc_hd__clkbuf_1 _08704_ (.A(_04530_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _08705_ (.A0(\fifo0.fifo_store[67][10] ),
    .A1(_04445_),
    .S(_04519_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _08706_ (.A(_04531_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _08707_ (.A0(\fifo0.fifo_store[67][11] ),
    .A1(_04447_),
    .S(_04519_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_1 _08708_ (.A(_04532_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _08709_ (.A0(\fifo0.fifo_store[67][12] ),
    .A1(_04494_),
    .S(_04519_),
    .X(_04533_));
 sky130_fd_sc_hd__clkbuf_1 _08710_ (.A(_04533_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _08711_ (.A0(\fifo0.fifo_store[67][13] ),
    .A1(_04468_),
    .S(_04519_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _08712_ (.A(_04534_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _08713_ (.A0(\fifo0.fifo_store[67][14] ),
    .A1(_04497_),
    .S(_04519_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _08714_ (.A(_04535_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _08715_ (.A0(\fifo0.fifo_store[67][15] ),
    .A1(_04499_),
    .S(_04519_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _08716_ (.A(_04536_),
    .X(_00518_));
 sky130_fd_sc_hd__nor2_4 _08717_ (.A(_03816_),
    .B(_04317_),
    .Y(_04537_));
 sky130_fd_sc_hd__buf_8 _08718_ (.A(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__mux2_1 _08719_ (.A0(\fifo0.fifo_store[112][0] ),
    .A1(_04472_),
    .S(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_1 _08720_ (.A(_04539_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _08721_ (.A0(\fifo0.fifo_store[112][1] ),
    .A1(_04476_),
    .S(_04538_),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_1 _08722_ (.A(_04540_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _08723_ (.A0(\fifo0.fifo_store[112][2] ),
    .A1(_04478_),
    .S(_04538_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_1 _08724_ (.A(_04541_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _08725_ (.A0(\fifo0.fifo_store[112][3] ),
    .A1(_04480_),
    .S(_04538_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _08726_ (.A(_04542_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _08727_ (.A0(\fifo0.fifo_store[112][4] ),
    .A1(_04482_),
    .S(_04538_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _08728_ (.A(_04543_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _08729_ (.A0(\fifo0.fifo_store[112][5] ),
    .A1(_04438_),
    .S(_04538_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _08730_ (.A(_04544_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _08731_ (.A0(\fifo0.fifo_store[112][6] ),
    .A1(_04485_),
    .S(_04538_),
    .X(_04545_));
 sky130_fd_sc_hd__clkbuf_1 _08732_ (.A(_04545_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _08733_ (.A0(\fifo0.fifo_store[112][7] ),
    .A1(_04441_),
    .S(_04538_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _08734_ (.A(_04546_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(\fifo0.fifo_store[112][8] ),
    .A1(_04488_),
    .S(_04538_),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_1 _08736_ (.A(_04547_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _08737_ (.A0(\fifo0.fifo_store[112][9] ),
    .A1(_04490_),
    .S(_04538_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _08738_ (.A(_04548_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _08739_ (.A0(\fifo0.fifo_store[112][10] ),
    .A1(_04445_),
    .S(_04537_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _08740_ (.A(_04549_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(\fifo0.fifo_store[112][11] ),
    .A1(_04447_),
    .S(_04537_),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _08742_ (.A(_04550_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _08743_ (.A0(\fifo0.fifo_store[112][12] ),
    .A1(_04494_),
    .S(_04537_),
    .X(_04551_));
 sky130_fd_sc_hd__clkbuf_1 _08744_ (.A(_04551_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _08745_ (.A0(\fifo0.fifo_store[112][13] ),
    .A1(_04468_),
    .S(_04537_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _08746_ (.A(_04552_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _08747_ (.A0(\fifo0.fifo_store[112][14] ),
    .A1(_04497_),
    .S(_04537_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_1 _08748_ (.A(_04553_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _08749_ (.A0(\fifo0.fifo_store[112][15] ),
    .A1(_04499_),
    .S(_04537_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _08750_ (.A(_04554_),
    .X(_00534_));
 sky130_fd_sc_hd__nor2_8 _08751_ (.A(_03986_),
    .B(_04277_),
    .Y(_04555_));
 sky130_fd_sc_hd__buf_6 _08752_ (.A(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_1 _08753_ (.A0(\fifo0.fifo_store[100][0] ),
    .A1(_04472_),
    .S(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _08754_ (.A(_04557_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(\fifo0.fifo_store[100][1] ),
    .A1(_04476_),
    .S(_04556_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _08756_ (.A(_04558_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _08757_ (.A0(\fifo0.fifo_store[100][2] ),
    .A1(_04478_),
    .S(_04556_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _08758_ (.A(_04559_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _08759_ (.A0(\fifo0.fifo_store[100][3] ),
    .A1(_04480_),
    .S(_04556_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _08760_ (.A(_04560_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _08761_ (.A0(\fifo0.fifo_store[100][4] ),
    .A1(_04482_),
    .S(_04556_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _08762_ (.A(_04561_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _08763_ (.A0(\fifo0.fifo_store[100][5] ),
    .A1(_04438_),
    .S(_04556_),
    .X(_04562_));
 sky130_fd_sc_hd__clkbuf_1 _08764_ (.A(_04562_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _08765_ (.A0(\fifo0.fifo_store[100][6] ),
    .A1(_04485_),
    .S(_04556_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _08766_ (.A(_04563_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _08767_ (.A0(\fifo0.fifo_store[100][7] ),
    .A1(_04441_),
    .S(_04556_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _08768_ (.A(_04564_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _08769_ (.A0(\fifo0.fifo_store[100][8] ),
    .A1(_04488_),
    .S(_04556_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _08770_ (.A(_04565_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _08771_ (.A0(\fifo0.fifo_store[100][9] ),
    .A1(_04490_),
    .S(_04556_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _08772_ (.A(_04566_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _08773_ (.A0(\fifo0.fifo_store[100][10] ),
    .A1(_04445_),
    .S(_04555_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _08774_ (.A(_04567_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _08775_ (.A0(\fifo0.fifo_store[100][11] ),
    .A1(_04447_),
    .S(_04555_),
    .X(_04568_));
 sky130_fd_sc_hd__clkbuf_1 _08776_ (.A(_04568_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _08777_ (.A0(\fifo0.fifo_store[100][12] ),
    .A1(_04494_),
    .S(_04555_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_1 _08778_ (.A(_04569_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _08779_ (.A0(\fifo0.fifo_store[100][13] ),
    .A1(_04468_),
    .S(_04555_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_1 _08780_ (.A(_04570_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _08781_ (.A0(\fifo0.fifo_store[100][14] ),
    .A1(_04497_),
    .S(_04555_),
    .X(_04571_));
 sky130_fd_sc_hd__clkbuf_1 _08782_ (.A(_04571_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _08783_ (.A0(\fifo0.fifo_store[100][15] ),
    .A1(_04499_),
    .S(_04555_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _08784_ (.A(_04572_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_4 _08785_ (.A(_04032_),
    .B(_04317_),
    .Y(_04573_));
 sky130_fd_sc_hd__buf_8 _08786_ (.A(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__mux2_1 _08787_ (.A0(\fifo0.fifo_store[113][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_1 _08788_ (.A(_04575_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _08789_ (.A0(\fifo0.fifo_store[113][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_04574_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _08790_ (.A(_04576_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _08791_ (.A0(\fifo0.fifo_store[113][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_04574_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _08792_ (.A(_04577_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(\fifo0.fifo_store[113][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_04574_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _08794_ (.A(_04578_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _08795_ (.A0(\fifo0.fifo_store[113][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_04574_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _08796_ (.A(_04579_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _08797_ (.A0(\fifo0.fifo_store[113][5] ),
    .A1(_04438_),
    .S(_04574_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _08798_ (.A(_04580_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _08799_ (.A0(\fifo0.fifo_store[113][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_04574_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_1 _08800_ (.A(_04581_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _08801_ (.A0(\fifo0.fifo_store[113][7] ),
    .A1(_04441_),
    .S(_04574_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _08802_ (.A(_04582_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _08803_ (.A0(\fifo0.fifo_store[113][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_04574_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _08804_ (.A(_04583_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(\fifo0.fifo_store[113][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_04574_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_1 _08806_ (.A(_04584_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(\fifo0.fifo_store[113][10] ),
    .A1(_04445_),
    .S(_04573_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _08808_ (.A(_04585_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(\fifo0.fifo_store[113][11] ),
    .A1(_04447_),
    .S(_04573_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _08810_ (.A(_04586_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(\fifo0.fifo_store[113][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_04573_),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_1 _08812_ (.A(_04587_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _08813_ (.A0(\fifo0.fifo_store[113][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_04573_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_1 _08814_ (.A(_04588_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(\fifo0.fifo_store[113][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_04573_),
    .X(_04589_));
 sky130_fd_sc_hd__clkbuf_1 _08816_ (.A(_04589_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _08817_ (.A0(\fifo0.fifo_store[113][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_04573_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _08818_ (.A(_04590_),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_8 _08819_ (.A(_03920_),
    .B(_04297_),
    .Y(_04591_));
 sky130_fd_sc_hd__buf_6 _08820_ (.A(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__mux2_1 _08821_ (.A0(\fifo0.fifo_store[111][0] ),
    .A1(_04472_),
    .S(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _08822_ (.A(_04593_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(\fifo0.fifo_store[111][1] ),
    .A1(_04476_),
    .S(_04592_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _08824_ (.A(_04594_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _08825_ (.A0(\fifo0.fifo_store[111][2] ),
    .A1(_04478_),
    .S(_04592_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _08826_ (.A(_04595_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _08827_ (.A0(\fifo0.fifo_store[111][3] ),
    .A1(_04480_),
    .S(_04592_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _08828_ (.A(_04596_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _08829_ (.A0(\fifo0.fifo_store[111][4] ),
    .A1(_04482_),
    .S(_04592_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _08830_ (.A(_04597_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _08831_ (.A0(\fifo0.fifo_store[111][5] ),
    .A1(_04438_),
    .S(_04592_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _08832_ (.A(_04598_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _08833_ (.A0(\fifo0.fifo_store[111][6] ),
    .A1(_04485_),
    .S(_04592_),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_1 _08834_ (.A(_04599_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _08835_ (.A0(\fifo0.fifo_store[111][7] ),
    .A1(_04441_),
    .S(_04592_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _08836_ (.A(_04600_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _08837_ (.A0(\fifo0.fifo_store[111][8] ),
    .A1(_04488_),
    .S(_04592_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _08838_ (.A(_04601_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(\fifo0.fifo_store[111][9] ),
    .A1(_04490_),
    .S(_04592_),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_1 _08840_ (.A(_04602_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(\fifo0.fifo_store[111][10] ),
    .A1(_04445_),
    .S(_04591_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_1 _08842_ (.A(_04603_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(\fifo0.fifo_store[111][11] ),
    .A1(_04447_),
    .S(_04591_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _08844_ (.A(_04604_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(\fifo0.fifo_store[111][12] ),
    .A1(_04494_),
    .S(_04591_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _08846_ (.A(_04605_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _08847_ (.A0(\fifo0.fifo_store[111][13] ),
    .A1(_04468_),
    .S(_04591_),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_1 _08848_ (.A(_04606_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _08849_ (.A0(\fifo0.fifo_store[111][14] ),
    .A1(_04497_),
    .S(_04591_),
    .X(_04607_));
 sky130_fd_sc_hd__clkbuf_1 _08850_ (.A(_04607_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _08851_ (.A0(\fifo0.fifo_store[111][15] ),
    .A1(_04499_),
    .S(_04591_),
    .X(_04608_));
 sky130_fd_sc_hd__clkbuf_1 _08852_ (.A(_04608_),
    .X(_00582_));
 sky130_fd_sc_hd__nor2_4 _08853_ (.A(_03990_),
    .B(_04317_),
    .Y(_04609_));
 sky130_fd_sc_hd__buf_8 _08854_ (.A(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__mux2_1 _08855_ (.A0(\fifo0.fifo_store[114][0] ),
    .A1(_04472_),
    .S(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__clkbuf_1 _08856_ (.A(_04611_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _08857_ (.A0(\fifo0.fifo_store[114][1] ),
    .A1(_04476_),
    .S(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _08858_ (.A(_04612_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _08859_ (.A0(\fifo0.fifo_store[114][2] ),
    .A1(_04478_),
    .S(_04610_),
    .X(_04613_));
 sky130_fd_sc_hd__clkbuf_1 _08860_ (.A(_04613_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _08861_ (.A0(\fifo0.fifo_store[114][3] ),
    .A1(_04480_),
    .S(_04610_),
    .X(_04614_));
 sky130_fd_sc_hd__clkbuf_1 _08862_ (.A(_04614_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _08863_ (.A0(\fifo0.fifo_store[114][4] ),
    .A1(_04482_),
    .S(_04610_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _08864_ (.A(_04615_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _08865_ (.A0(\fifo0.fifo_store[114][5] ),
    .A1(_04438_),
    .S(_04610_),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_1 _08866_ (.A(_04616_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _08867_ (.A0(\fifo0.fifo_store[114][6] ),
    .A1(_04485_),
    .S(_04610_),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_1 _08868_ (.A(_04617_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _08869_ (.A0(\fifo0.fifo_store[114][7] ),
    .A1(_04441_),
    .S(_04610_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_1 _08870_ (.A(_04618_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _08871_ (.A0(\fifo0.fifo_store[114][8] ),
    .A1(_04488_),
    .S(_04610_),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _08872_ (.A(_04619_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _08873_ (.A0(\fifo0.fifo_store[114][9] ),
    .A1(_04490_),
    .S(_04610_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _08874_ (.A(_04620_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(\fifo0.fifo_store[114][10] ),
    .A1(_04445_),
    .S(_04609_),
    .X(_04621_));
 sky130_fd_sc_hd__clkbuf_1 _08876_ (.A(_04621_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _08877_ (.A0(\fifo0.fifo_store[114][11] ),
    .A1(_04447_),
    .S(_04609_),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_1 _08878_ (.A(_04622_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(\fifo0.fifo_store[114][12] ),
    .A1(_04494_),
    .S(_04609_),
    .X(_04623_));
 sky130_fd_sc_hd__clkbuf_1 _08880_ (.A(_04623_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _08881_ (.A0(\fifo0.fifo_store[114][13] ),
    .A1(_04468_),
    .S(_04609_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _08882_ (.A(_04624_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(\fifo0.fifo_store[114][14] ),
    .A1(_04497_),
    .S(_04609_),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _08884_ (.A(_04625_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(\fifo0.fifo_store[114][15] ),
    .A1(_04499_),
    .S(_04609_),
    .X(_04626_));
 sky130_fd_sc_hd__clkbuf_1 _08886_ (.A(_04626_),
    .X(_00598_));
 sky130_fd_sc_hd__nand2_2 _08887_ (.A(_03810_),
    .B(_03809_),
    .Y(_04627_));
 sky130_fd_sc_hd__or2_1 _08888_ (.A(_03939_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__buf_12 _08889_ (.A(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__or2_1 _08890_ (.A(_04201_),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__buf_6 _08891_ (.A(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__buf_8 _08892_ (.A(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__mux2_1 _08893_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[46][0] ),
    .S(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _08894_ (.A(_04633_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _08895_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[46][1] ),
    .S(_04632_),
    .X(_04634_));
 sky130_fd_sc_hd__clkbuf_1 _08896_ (.A(_04634_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _08897_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[46][2] ),
    .S(_04632_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _08898_ (.A(_04635_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[46][3] ),
    .S(_04632_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _08900_ (.A(_04636_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _08901_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[46][4] ),
    .S(_04632_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _08902_ (.A(_04637_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _08903_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[46][5] ),
    .S(_04632_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _08904_ (.A(_04638_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _08905_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[46][6] ),
    .S(_04632_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _08906_ (.A(_04639_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _08907_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[46][7] ),
    .S(_04632_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_1 _08908_ (.A(_04640_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _08909_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[46][8] ),
    .S(_04632_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _08910_ (.A(_04641_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _08911_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[46][9] ),
    .S(_04632_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _08912_ (.A(_04642_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _08913_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[46][10] ),
    .S(_04631_),
    .X(_04643_));
 sky130_fd_sc_hd__clkbuf_1 _08914_ (.A(_04643_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _08915_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[46][11] ),
    .S(_04631_),
    .X(_04644_));
 sky130_fd_sc_hd__clkbuf_1 _08916_ (.A(_04644_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _08917_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[46][12] ),
    .S(_04631_),
    .X(_04645_));
 sky130_fd_sc_hd__clkbuf_1 _08918_ (.A(_04645_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _08919_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[46][13] ),
    .S(_04631_),
    .X(_04646_));
 sky130_fd_sc_hd__clkbuf_1 _08920_ (.A(_04646_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _08921_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[46][14] ),
    .S(_04631_),
    .X(_04647_));
 sky130_fd_sc_hd__clkbuf_1 _08922_ (.A(_04647_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[46][15] ),
    .S(_04631_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_1 _08924_ (.A(_04648_),
    .X(_00614_));
 sky130_fd_sc_hd__nor2_8 _08925_ (.A(_04053_),
    .B(_04172_),
    .Y(_04649_));
 sky130_fd_sc_hd__buf_12 _08926_ (.A(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(\fifo0.fifo_store[91][0] ),
    .A1(_04472_),
    .S(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_1 _08928_ (.A(_04651_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _08929_ (.A0(\fifo0.fifo_store[91][1] ),
    .A1(_04476_),
    .S(_04650_),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_1 _08930_ (.A(_04652_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(\fifo0.fifo_store[91][2] ),
    .A1(_04478_),
    .S(_04650_),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_1 _08932_ (.A(_04653_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(\fifo0.fifo_store[91][3] ),
    .A1(_04480_),
    .S(_04650_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_1 _08934_ (.A(_04654_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _08935_ (.A0(\fifo0.fifo_store[91][4] ),
    .A1(_04482_),
    .S(_04650_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_1 _08936_ (.A(_04655_),
    .X(_00619_));
 sky130_fd_sc_hd__buf_4 _08937_ (.A(_03838_),
    .X(_04656_));
 sky130_fd_sc_hd__mux2_1 _08938_ (.A0(\fifo0.fifo_store[91][5] ),
    .A1(_04656_),
    .S(_04650_),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_1 _08939_ (.A(_04657_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(\fifo0.fifo_store[91][6] ),
    .A1(_04485_),
    .S(_04650_),
    .X(_04658_));
 sky130_fd_sc_hd__clkbuf_1 _08941_ (.A(_04658_),
    .X(_00621_));
 sky130_fd_sc_hd__clkbuf_4 _08942_ (.A(_03843_),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_1 _08943_ (.A0(\fifo0.fifo_store[91][7] ),
    .A1(_04659_),
    .S(_04650_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _08944_ (.A(_04660_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(\fifo0.fifo_store[91][8] ),
    .A1(_04488_),
    .S(_04650_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _08946_ (.A(_04661_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(\fifo0.fifo_store[91][9] ),
    .A1(_04490_),
    .S(_04650_),
    .X(_04662_));
 sky130_fd_sc_hd__clkbuf_1 _08948_ (.A(_04662_),
    .X(_00624_));
 sky130_fd_sc_hd__buf_4 _08949_ (.A(_03850_),
    .X(_04663_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(\fifo0.fifo_store[91][10] ),
    .A1(_04663_),
    .S(_04649_),
    .X(_04664_));
 sky130_fd_sc_hd__clkbuf_1 _08951_ (.A(_04664_),
    .X(_00625_));
 sky130_fd_sc_hd__buf_4 _08952_ (.A(_03853_),
    .X(_04665_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(\fifo0.fifo_store[91][11] ),
    .A1(_04665_),
    .S(_04649_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _08954_ (.A(_04666_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(\fifo0.fifo_store[91][12] ),
    .A1(_04494_),
    .S(_04649_),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _08956_ (.A(_04667_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _08957_ (.A0(\fifo0.fifo_store[91][13] ),
    .A1(_04468_),
    .S(_04649_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_1 _08958_ (.A(_04668_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(\fifo0.fifo_store[91][14] ),
    .A1(_04497_),
    .S(_04649_),
    .X(_04669_));
 sky130_fd_sc_hd__clkbuf_1 _08960_ (.A(_04669_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _08961_ (.A0(\fifo0.fifo_store[91][15] ),
    .A1(_04499_),
    .S(_04649_),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_1 _08962_ (.A(_04670_),
    .X(_00630_));
 sky130_fd_sc_hd__nor2_4 _08963_ (.A(_03990_),
    .B(_04145_),
    .Y(_04671_));
 sky130_fd_sc_hd__buf_6 _08964_ (.A(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _08965_ (.A0(\fifo0.fifo_store[66][0] ),
    .A1(_04472_),
    .S(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _08966_ (.A(_04673_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(\fifo0.fifo_store[66][1] ),
    .A1(_04476_),
    .S(_04672_),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_1 _08968_ (.A(_04674_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(\fifo0.fifo_store[66][2] ),
    .A1(_04478_),
    .S(_04672_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _08970_ (.A(_04675_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(\fifo0.fifo_store[66][3] ),
    .A1(_04480_),
    .S(_04672_),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_1 _08972_ (.A(_04676_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(\fifo0.fifo_store[66][4] ),
    .A1(_04482_),
    .S(_04672_),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _08974_ (.A(_04677_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(\fifo0.fifo_store[66][5] ),
    .A1(_04656_),
    .S(_04672_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _08976_ (.A(_04678_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _08977_ (.A0(\fifo0.fifo_store[66][6] ),
    .A1(_04485_),
    .S(_04672_),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _08978_ (.A(_04679_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(\fifo0.fifo_store[66][7] ),
    .A1(_04659_),
    .S(_04672_),
    .X(_04680_));
 sky130_fd_sc_hd__clkbuf_1 _08980_ (.A(_04680_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _08981_ (.A0(\fifo0.fifo_store[66][8] ),
    .A1(_04488_),
    .S(_04672_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _08982_ (.A(_04681_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(\fifo0.fifo_store[66][9] ),
    .A1(_04490_),
    .S(_04672_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_1 _08984_ (.A(_04682_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _08985_ (.A0(\fifo0.fifo_store[66][10] ),
    .A1(_04663_),
    .S(_04671_),
    .X(_04683_));
 sky130_fd_sc_hd__clkbuf_1 _08986_ (.A(_04683_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(\fifo0.fifo_store[66][11] ),
    .A1(_04665_),
    .S(_04671_),
    .X(_04684_));
 sky130_fd_sc_hd__clkbuf_1 _08988_ (.A(_04684_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _08989_ (.A0(\fifo0.fifo_store[66][12] ),
    .A1(_04494_),
    .S(_04671_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_1 _08990_ (.A(_04685_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _08991_ (.A0(\fifo0.fifo_store[66][13] ),
    .A1(_04468_),
    .S(_04671_),
    .X(_04686_));
 sky130_fd_sc_hd__clkbuf_1 _08992_ (.A(_04686_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(\fifo0.fifo_store[66][14] ),
    .A1(_04497_),
    .S(_04671_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _08994_ (.A(_04687_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(\fifo0.fifo_store[66][15] ),
    .A1(_04499_),
    .S(_04671_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _08996_ (.A(_04688_),
    .X(_00646_));
 sky130_fd_sc_hd__or2_1 _08997_ (.A(_03865_),
    .B(_04627_),
    .X(_04689_));
 sky130_fd_sc_hd__buf_12 _08998_ (.A(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__nor2_8 _08999_ (.A(_04032_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__buf_6 _09000_ (.A(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_1 _09001_ (.A0(\fifo0.fifo_store[49][0] ),
    .A1(_04472_),
    .S(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _09002_ (.A(_04693_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(\fifo0.fifo_store[49][1] ),
    .A1(_04476_),
    .S(_04692_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _09004_ (.A(_04694_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(\fifo0.fifo_store[49][2] ),
    .A1(_04478_),
    .S(_04692_),
    .X(_04695_));
 sky130_fd_sc_hd__clkbuf_1 _09006_ (.A(_04695_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _09007_ (.A0(\fifo0.fifo_store[49][3] ),
    .A1(_04480_),
    .S(_04692_),
    .X(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _09008_ (.A(_04696_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _09009_ (.A0(\fifo0.fifo_store[49][4] ),
    .A1(_04482_),
    .S(_04692_),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_1 _09010_ (.A(_04697_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(\fifo0.fifo_store[49][5] ),
    .A1(_04656_),
    .S(_04692_),
    .X(_04698_));
 sky130_fd_sc_hd__clkbuf_1 _09012_ (.A(_04698_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _09013_ (.A0(\fifo0.fifo_store[49][6] ),
    .A1(_04485_),
    .S(_04692_),
    .X(_04699_));
 sky130_fd_sc_hd__clkbuf_1 _09014_ (.A(_04699_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _09015_ (.A0(\fifo0.fifo_store[49][7] ),
    .A1(_04659_),
    .S(_04692_),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_1 _09016_ (.A(_04700_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _09017_ (.A0(\fifo0.fifo_store[49][8] ),
    .A1(_04488_),
    .S(_04692_),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _09018_ (.A(_04701_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _09019_ (.A0(\fifo0.fifo_store[49][9] ),
    .A1(_04490_),
    .S(_04692_),
    .X(_04702_));
 sky130_fd_sc_hd__clkbuf_1 _09020_ (.A(_04702_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(\fifo0.fifo_store[49][10] ),
    .A1(_04663_),
    .S(_04691_),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_1 _09022_ (.A(_04703_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(\fifo0.fifo_store[49][11] ),
    .A1(_04665_),
    .S(_04691_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_1 _09024_ (.A(_04704_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _09025_ (.A0(\fifo0.fifo_store[49][12] ),
    .A1(_04494_),
    .S(_04691_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _09026_ (.A(_04705_),
    .X(_00659_));
 sky130_fd_sc_hd__buf_6 _09027_ (.A(_03908_),
    .X(_04706_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(\fifo0.fifo_store[49][13] ),
    .A1(_04706_),
    .S(_04691_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _09029_ (.A(_04707_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _09030_ (.A0(\fifo0.fifo_store[49][14] ),
    .A1(_04497_),
    .S(_04691_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _09031_ (.A(_04708_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(\fifo0.fifo_store[49][15] ),
    .A1(_04499_),
    .S(_04691_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _09033_ (.A(_04709_),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _09034_ (.A(_04201_),
    .B(_04297_),
    .X(_04710_));
 sky130_fd_sc_hd__buf_4 _09035_ (.A(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__buf_6 _09036_ (.A(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__mux2_1 _09037_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[110][0] ),
    .S(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _09038_ (.A(_04713_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[110][1] ),
    .S(_04712_),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _09040_ (.A(_04714_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[110][2] ),
    .S(_04712_),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_1 _09042_ (.A(_04715_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[110][3] ),
    .S(_04712_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_1 _09044_ (.A(_04716_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[110][4] ),
    .S(_04712_),
    .X(_04717_));
 sky130_fd_sc_hd__clkbuf_1 _09046_ (.A(_04717_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[110][5] ),
    .S(_04712_),
    .X(_04718_));
 sky130_fd_sc_hd__clkbuf_1 _09048_ (.A(_04718_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[110][6] ),
    .S(_04712_),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_1 _09050_ (.A(_04719_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[110][7] ),
    .S(_04712_),
    .X(_04720_));
 sky130_fd_sc_hd__clkbuf_1 _09052_ (.A(_04720_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _09053_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[110][8] ),
    .S(_04712_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _09054_ (.A(_04721_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _09055_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[110][9] ),
    .S(_04712_),
    .X(_04722_));
 sky130_fd_sc_hd__clkbuf_1 _09056_ (.A(_04722_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _09057_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[110][10] ),
    .S(_04711_),
    .X(_04723_));
 sky130_fd_sc_hd__clkbuf_1 _09058_ (.A(_04723_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[110][11] ),
    .S(_04711_),
    .X(_04724_));
 sky130_fd_sc_hd__clkbuf_1 _09060_ (.A(_04724_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _09061_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[110][12] ),
    .S(_04711_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _09062_ (.A(_04725_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[110][13] ),
    .S(_04711_),
    .X(_04726_));
 sky130_fd_sc_hd__clkbuf_1 _09064_ (.A(_04726_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _09065_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[110][14] ),
    .S(_04711_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _09066_ (.A(_04727_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _09067_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[110][15] ),
    .S(_04711_),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_1 _09068_ (.A(_04728_),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_4 _09069_ (.A(_03821_),
    .X(_04729_));
 sky130_fd_sc_hd__nor2_8 _09070_ (.A(_03816_),
    .B(_04297_),
    .Y(_04730_));
 sky130_fd_sc_hd__buf_12 _09071_ (.A(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(\fifo0.fifo_store[104][0] ),
    .A1(_04729_),
    .S(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__clkbuf_1 _09073_ (.A(_04732_),
    .X(_00679_));
 sky130_fd_sc_hd__buf_4 _09074_ (.A(_03872_),
    .X(_04733_));
 sky130_fd_sc_hd__mux2_1 _09075_ (.A0(\fifo0.fifo_store[104][1] ),
    .A1(_04733_),
    .S(_04731_),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_1 _09076_ (.A(_04734_),
    .X(_00680_));
 sky130_fd_sc_hd__buf_4 _09077_ (.A(_03875_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(\fifo0.fifo_store[104][2] ),
    .A1(_04735_),
    .S(_04731_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _09079_ (.A(_04736_),
    .X(_00681_));
 sky130_fd_sc_hd__buf_4 _09080_ (.A(_03878_),
    .X(_04737_));
 sky130_fd_sc_hd__mux2_1 _09081_ (.A0(\fifo0.fifo_store[104][3] ),
    .A1(_04737_),
    .S(_04731_),
    .X(_04738_));
 sky130_fd_sc_hd__clkbuf_1 _09082_ (.A(_04738_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_4 _09083_ (.A(_03881_),
    .X(_04739_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(\fifo0.fifo_store[104][4] ),
    .A1(_04739_),
    .S(_04731_),
    .X(_04740_));
 sky130_fd_sc_hd__clkbuf_1 _09085_ (.A(_04740_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(\fifo0.fifo_store[104][5] ),
    .A1(_04656_),
    .S(_04731_),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_1 _09087_ (.A(_04741_),
    .X(_00684_));
 sky130_fd_sc_hd__buf_4 _09088_ (.A(_03887_),
    .X(_04742_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(\fifo0.fifo_store[104][6] ),
    .A1(_04742_),
    .S(_04731_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _09090_ (.A(_04743_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _09091_ (.A0(\fifo0.fifo_store[104][7] ),
    .A1(_04659_),
    .S(_04731_),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_1 _09092_ (.A(_04744_),
    .X(_00686_));
 sky130_fd_sc_hd__buf_4 _09093_ (.A(_03893_),
    .X(_04745_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(\fifo0.fifo_store[104][8] ),
    .A1(_04745_),
    .S(_04731_),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_1 _09095_ (.A(_04746_),
    .X(_00687_));
 sky130_fd_sc_hd__clkbuf_4 _09096_ (.A(_03896_),
    .X(_04747_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(\fifo0.fifo_store[104][9] ),
    .A1(_04747_),
    .S(_04731_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _09098_ (.A(_04748_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(\fifo0.fifo_store[104][10] ),
    .A1(_04663_),
    .S(_04730_),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_1 _09100_ (.A(_04749_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _09101_ (.A0(\fifo0.fifo_store[104][11] ),
    .A1(_04665_),
    .S(_04730_),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_1 _09102_ (.A(_04750_),
    .X(_00690_));
 sky130_fd_sc_hd__buf_4 _09103_ (.A(_03905_),
    .X(_04751_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(\fifo0.fifo_store[104][12] ),
    .A1(_04751_),
    .S(_04730_),
    .X(_04752_));
 sky130_fd_sc_hd__clkbuf_1 _09105_ (.A(_04752_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(\fifo0.fifo_store[104][13] ),
    .A1(_04706_),
    .S(_04730_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_1 _09107_ (.A(_04753_),
    .X(_00692_));
 sky130_fd_sc_hd__buf_4 _09108_ (.A(_03911_),
    .X(_04754_));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(\fifo0.fifo_store[104][14] ),
    .A1(_04754_),
    .S(_04730_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_1 _09110_ (.A(_04755_),
    .X(_00693_));
 sky130_fd_sc_hd__buf_4 _09111_ (.A(_03914_),
    .X(_04756_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(\fifo0.fifo_store[104][15] ),
    .A1(_04756_),
    .S(_04730_),
    .X(_04757_));
 sky130_fd_sc_hd__clkbuf_1 _09113_ (.A(_04757_),
    .X(_00694_));
 sky130_fd_sc_hd__nor2_8 _09114_ (.A(_03990_),
    .B(_04356_),
    .Y(_04758_));
 sky130_fd_sc_hd__buf_12 _09115_ (.A(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(\fifo0.fifo_store[10][0] ),
    .A1(_04729_),
    .S(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__clkbuf_1 _09117_ (.A(_04760_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(\fifo0.fifo_store[10][1] ),
    .A1(_04733_),
    .S(_04759_),
    .X(_04761_));
 sky130_fd_sc_hd__clkbuf_1 _09119_ (.A(_04761_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(\fifo0.fifo_store[10][2] ),
    .A1(_04735_),
    .S(_04759_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_1 _09121_ (.A(_04762_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(\fifo0.fifo_store[10][3] ),
    .A1(_04737_),
    .S(_04759_),
    .X(_04763_));
 sky130_fd_sc_hd__clkbuf_1 _09123_ (.A(_04763_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(\fifo0.fifo_store[10][4] ),
    .A1(_04739_),
    .S(_04759_),
    .X(_04764_));
 sky130_fd_sc_hd__clkbuf_1 _09125_ (.A(_04764_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(\fifo0.fifo_store[10][5] ),
    .A1(_04656_),
    .S(_04759_),
    .X(_04765_));
 sky130_fd_sc_hd__clkbuf_1 _09127_ (.A(_04765_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(\fifo0.fifo_store[10][6] ),
    .A1(_04742_),
    .S(_04759_),
    .X(_04766_));
 sky130_fd_sc_hd__clkbuf_1 _09129_ (.A(_04766_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(\fifo0.fifo_store[10][7] ),
    .A1(_04659_),
    .S(_04759_),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_1 _09131_ (.A(_04767_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(\fifo0.fifo_store[10][8] ),
    .A1(_04745_),
    .S(_04759_),
    .X(_04768_));
 sky130_fd_sc_hd__clkbuf_1 _09133_ (.A(_04768_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(\fifo0.fifo_store[10][9] ),
    .A1(_04747_),
    .S(_04759_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_1 _09135_ (.A(_04769_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(\fifo0.fifo_store[10][10] ),
    .A1(_04663_),
    .S(_04758_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_1 _09137_ (.A(_04770_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(\fifo0.fifo_store[10][11] ),
    .A1(_04665_),
    .S(_04758_),
    .X(_04771_));
 sky130_fd_sc_hd__clkbuf_1 _09139_ (.A(_04771_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(\fifo0.fifo_store[10][12] ),
    .A1(_04751_),
    .S(_04758_),
    .X(_04772_));
 sky130_fd_sc_hd__clkbuf_1 _09141_ (.A(_04772_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(\fifo0.fifo_store[10][13] ),
    .A1(_04706_),
    .S(_04758_),
    .X(_04773_));
 sky130_fd_sc_hd__clkbuf_1 _09143_ (.A(_04773_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(\fifo0.fifo_store[10][14] ),
    .A1(_04754_),
    .S(_04758_),
    .X(_04774_));
 sky130_fd_sc_hd__clkbuf_1 _09145_ (.A(_04774_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(\fifo0.fifo_store[10][15] ),
    .A1(_04756_),
    .S(_04758_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_1 _09147_ (.A(_04775_),
    .X(_00710_));
 sky130_fd_sc_hd__nor2_8 _09148_ (.A(_03920_),
    .B(_03986_),
    .Y(_04776_));
 sky130_fd_sc_hd__buf_8 _09149_ (.A(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(\fifo0.fifo_store[103][0] ),
    .A1(_04729_),
    .S(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__clkbuf_1 _09151_ (.A(_04778_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _09152_ (.A0(\fifo0.fifo_store[103][1] ),
    .A1(_04733_),
    .S(_04777_),
    .X(_04779_));
 sky130_fd_sc_hd__clkbuf_1 _09153_ (.A(_04779_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(\fifo0.fifo_store[103][2] ),
    .A1(_04735_),
    .S(_04777_),
    .X(_04780_));
 sky130_fd_sc_hd__clkbuf_1 _09155_ (.A(_04780_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(\fifo0.fifo_store[103][3] ),
    .A1(_04737_),
    .S(_04777_),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_1 _09157_ (.A(_04781_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(\fifo0.fifo_store[103][4] ),
    .A1(_04739_),
    .S(_04777_),
    .X(_04782_));
 sky130_fd_sc_hd__clkbuf_1 _09159_ (.A(_04782_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(\fifo0.fifo_store[103][5] ),
    .A1(_04656_),
    .S(_04777_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_1 _09161_ (.A(_04783_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(\fifo0.fifo_store[103][6] ),
    .A1(_04742_),
    .S(_04777_),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_1 _09163_ (.A(_04784_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(\fifo0.fifo_store[103][7] ),
    .A1(_04659_),
    .S(_04777_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_1 _09165_ (.A(_04785_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(\fifo0.fifo_store[103][8] ),
    .A1(_04745_),
    .S(_04777_),
    .X(_04786_));
 sky130_fd_sc_hd__clkbuf_1 _09167_ (.A(_04786_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(\fifo0.fifo_store[103][9] ),
    .A1(_04747_),
    .S(_04777_),
    .X(_04787_));
 sky130_fd_sc_hd__clkbuf_1 _09169_ (.A(_04787_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(\fifo0.fifo_store[103][10] ),
    .A1(_04663_),
    .S(_04776_),
    .X(_04788_));
 sky130_fd_sc_hd__clkbuf_1 _09171_ (.A(_04788_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(\fifo0.fifo_store[103][11] ),
    .A1(_04665_),
    .S(_04776_),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_1 _09173_ (.A(_04789_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(\fifo0.fifo_store[103][12] ),
    .A1(_04751_),
    .S(_04776_),
    .X(_04790_));
 sky130_fd_sc_hd__clkbuf_1 _09175_ (.A(_04790_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(\fifo0.fifo_store[103][13] ),
    .A1(_04706_),
    .S(_04776_),
    .X(_04791_));
 sky130_fd_sc_hd__clkbuf_1 _09177_ (.A(_04791_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(\fifo0.fifo_store[103][14] ),
    .A1(_04754_),
    .S(_04776_),
    .X(_04792_));
 sky130_fd_sc_hd__clkbuf_1 _09179_ (.A(_04792_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(\fifo0.fifo_store[103][15] ),
    .A1(_04756_),
    .S(_04776_),
    .X(_04793_));
 sky130_fd_sc_hd__clkbuf_1 _09181_ (.A(_04793_),
    .X(_00726_));
 sky130_fd_sc_hd__nor2_8 _09182_ (.A(_04277_),
    .B(_04297_),
    .Y(_04794_));
 sky130_fd_sc_hd__buf_6 _09183_ (.A(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(\fifo0.fifo_store[108][0] ),
    .A1(_04729_),
    .S(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__clkbuf_1 _09185_ (.A(_04796_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(\fifo0.fifo_store[108][1] ),
    .A1(_04733_),
    .S(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__clkbuf_1 _09187_ (.A(_04797_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(\fifo0.fifo_store[108][2] ),
    .A1(_04735_),
    .S(_04795_),
    .X(_04798_));
 sky130_fd_sc_hd__clkbuf_1 _09189_ (.A(_04798_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(\fifo0.fifo_store[108][3] ),
    .A1(_04737_),
    .S(_04795_),
    .X(_04799_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_04799_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(\fifo0.fifo_store[108][4] ),
    .A1(_04739_),
    .S(_04795_),
    .X(_04800_));
 sky130_fd_sc_hd__clkbuf_1 _09193_ (.A(_04800_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(\fifo0.fifo_store[108][5] ),
    .A1(_04656_),
    .S(_04795_),
    .X(_04801_));
 sky130_fd_sc_hd__clkbuf_1 _09195_ (.A(_04801_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(\fifo0.fifo_store[108][6] ),
    .A1(_04742_),
    .S(_04795_),
    .X(_04802_));
 sky130_fd_sc_hd__clkbuf_1 _09197_ (.A(_04802_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(\fifo0.fifo_store[108][7] ),
    .A1(_04659_),
    .S(_04795_),
    .X(_04803_));
 sky130_fd_sc_hd__clkbuf_1 _09199_ (.A(_04803_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(\fifo0.fifo_store[108][8] ),
    .A1(_04745_),
    .S(_04795_),
    .X(_04804_));
 sky130_fd_sc_hd__clkbuf_1 _09201_ (.A(_04804_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(\fifo0.fifo_store[108][9] ),
    .A1(_04747_),
    .S(_04795_),
    .X(_04805_));
 sky130_fd_sc_hd__clkbuf_1 _09203_ (.A(_04805_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(\fifo0.fifo_store[108][10] ),
    .A1(_04663_),
    .S(_04794_),
    .X(_04806_));
 sky130_fd_sc_hd__clkbuf_1 _09205_ (.A(_04806_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(\fifo0.fifo_store[108][11] ),
    .A1(_04665_),
    .S(_04794_),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_1 _09207_ (.A(_04807_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(\fifo0.fifo_store[108][12] ),
    .A1(_04751_),
    .S(_04794_),
    .X(_04808_));
 sky130_fd_sc_hd__clkbuf_1 _09209_ (.A(_04808_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(\fifo0.fifo_store[108][13] ),
    .A1(_04706_),
    .S(_04794_),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_1 _09211_ (.A(_04809_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(\fifo0.fifo_store[108][14] ),
    .A1(_04754_),
    .S(_04794_),
    .X(_04810_));
 sky130_fd_sc_hd__clkbuf_1 _09213_ (.A(_04810_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(\fifo0.fifo_store[108][15] ),
    .A1(_04756_),
    .S(_04794_),
    .X(_04811_));
 sky130_fd_sc_hd__clkbuf_1 _09215_ (.A(_04811_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _09216_ (.A(_04201_),
    .B(_03986_),
    .X(_04812_));
 sky130_fd_sc_hd__buf_4 _09217_ (.A(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__buf_6 _09218_ (.A(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(_03822_),
    .A1(\fifo0.fifo_store[102][0] ),
    .S(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__clkbuf_1 _09220_ (.A(_04815_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(_03829_),
    .A1(\fifo0.fifo_store[102][1] ),
    .S(_04814_),
    .X(_04816_));
 sky130_fd_sc_hd__clkbuf_1 _09222_ (.A(_04816_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(_03832_),
    .A1(\fifo0.fifo_store[102][2] ),
    .S(_04814_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _09224_ (.A(_04817_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(_03834_),
    .A1(\fifo0.fifo_store[102][3] ),
    .S(_04814_),
    .X(_04818_));
 sky130_fd_sc_hd__clkbuf_1 _09226_ (.A(_04818_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(_03836_),
    .A1(\fifo0.fifo_store[102][4] ),
    .S(_04814_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _09228_ (.A(_04819_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(_03839_),
    .A1(\fifo0.fifo_store[102][5] ),
    .S(_04814_),
    .X(_04820_));
 sky130_fd_sc_hd__clkbuf_1 _09230_ (.A(_04820_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(_03841_),
    .A1(\fifo0.fifo_store[102][6] ),
    .S(_04814_),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_1 _09232_ (.A(_04821_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(_03844_),
    .A1(\fifo0.fifo_store[102][7] ),
    .S(_04814_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_1 _09234_ (.A(_04822_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(_03846_),
    .A1(\fifo0.fifo_store[102][8] ),
    .S(_04814_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_1 _09236_ (.A(_04823_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(_03848_),
    .A1(\fifo0.fifo_store[102][9] ),
    .S(_04814_),
    .X(_04824_));
 sky130_fd_sc_hd__clkbuf_1 _09238_ (.A(_04824_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _09239_ (.A0(_03851_),
    .A1(\fifo0.fifo_store[102][10] ),
    .S(_04813_),
    .X(_04825_));
 sky130_fd_sc_hd__clkbuf_1 _09240_ (.A(_04825_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _09241_ (.A0(_03854_),
    .A1(\fifo0.fifo_store[102][11] ),
    .S(_04813_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_1 _09242_ (.A(_04826_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(_03856_),
    .A1(\fifo0.fifo_store[102][12] ),
    .S(_04813_),
    .X(_04827_));
 sky130_fd_sc_hd__clkbuf_1 _09244_ (.A(_04827_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _09245_ (.A0(_03858_),
    .A1(\fifo0.fifo_store[102][13] ),
    .S(_04813_),
    .X(_04828_));
 sky130_fd_sc_hd__clkbuf_1 _09246_ (.A(_04828_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(_03860_),
    .A1(\fifo0.fifo_store[102][14] ),
    .S(_04813_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _09248_ (.A(_04829_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(_03862_),
    .A1(\fifo0.fifo_store[102][15] ),
    .S(_04813_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_1 _09250_ (.A(_04830_),
    .X(_00758_));
 sky130_fd_sc_hd__nor2_8 _09251_ (.A(_03965_),
    .B(_03986_),
    .Y(_04831_));
 sky130_fd_sc_hd__buf_8 _09252_ (.A(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(\fifo0.fifo_store[101][0] ),
    .A1(_04729_),
    .S(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _09254_ (.A(_04833_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(\fifo0.fifo_store[101][1] ),
    .A1(_04733_),
    .S(_04832_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_1 _09256_ (.A(_04834_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(\fifo0.fifo_store[101][2] ),
    .A1(_04735_),
    .S(_04832_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _09258_ (.A(_04835_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(\fifo0.fifo_store[101][3] ),
    .A1(_04737_),
    .S(_04832_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _09260_ (.A(_04836_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _09261_ (.A0(\fifo0.fifo_store[101][4] ),
    .A1(_04739_),
    .S(_04832_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _09262_ (.A(_04837_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(\fifo0.fifo_store[101][5] ),
    .A1(_04656_),
    .S(_04832_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_1 _09264_ (.A(_04838_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(\fifo0.fifo_store[101][6] ),
    .A1(_04742_),
    .S(_04832_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _09266_ (.A(_04839_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(\fifo0.fifo_store[101][7] ),
    .A1(_04659_),
    .S(_04832_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _09268_ (.A(_04840_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(\fifo0.fifo_store[101][8] ),
    .A1(_04745_),
    .S(_04832_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _09270_ (.A(_04841_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _09271_ (.A0(\fifo0.fifo_store[101][9] ),
    .A1(_04747_),
    .S(_04832_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _09272_ (.A(_04842_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(\fifo0.fifo_store[101][10] ),
    .A1(_04663_),
    .S(_04831_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _09274_ (.A(_04843_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _09275_ (.A0(\fifo0.fifo_store[101][11] ),
    .A1(_04665_),
    .S(_04831_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _09276_ (.A(_04844_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(\fifo0.fifo_store[101][12] ),
    .A1(_04751_),
    .S(_04831_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _09278_ (.A(_04845_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(\fifo0.fifo_store[101][13] ),
    .A1(_04706_),
    .S(_04831_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _09280_ (.A(_04846_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(\fifo0.fifo_store[101][14] ),
    .A1(_04754_),
    .S(_04831_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _09282_ (.A(_04847_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(\fifo0.fifo_store[101][15] ),
    .A1(_04756_),
    .S(_04831_),
    .X(_04848_));
 sky130_fd_sc_hd__clkbuf_1 _09284_ (.A(_04848_),
    .X(_00774_));
 sky130_fd_sc_hd__nor2_8 _09285_ (.A(_04053_),
    .B(_04297_),
    .Y(_04849_));
 sky130_fd_sc_hd__clkbuf_16 _09286_ (.A(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(\fifo0.fifo_store[107][0] ),
    .A1(_04729_),
    .S(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_1 _09288_ (.A(_04851_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(\fifo0.fifo_store[107][1] ),
    .A1(_04733_),
    .S(_04850_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _09290_ (.A(_04852_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(\fifo0.fifo_store[107][2] ),
    .A1(_04735_),
    .S(_04850_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _09292_ (.A(_04853_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(\fifo0.fifo_store[107][3] ),
    .A1(_04737_),
    .S(_04850_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _09294_ (.A(_04854_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(\fifo0.fifo_store[107][4] ),
    .A1(_04739_),
    .S(_04850_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _09296_ (.A(_04855_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(\fifo0.fifo_store[107][5] ),
    .A1(_04656_),
    .S(_04850_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_1 _09298_ (.A(_04856_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(\fifo0.fifo_store[107][6] ),
    .A1(_04742_),
    .S(_04850_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _09300_ (.A(_04857_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(\fifo0.fifo_store[107][7] ),
    .A1(_04659_),
    .S(_04850_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _09302_ (.A(_04858_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(\fifo0.fifo_store[107][8] ),
    .A1(_04745_),
    .S(_04850_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _09304_ (.A(_04859_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(\fifo0.fifo_store[107][9] ),
    .A1(_04747_),
    .S(_04850_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _09306_ (.A(_04860_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(\fifo0.fifo_store[107][10] ),
    .A1(_04663_),
    .S(_04849_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _09308_ (.A(_04861_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(\fifo0.fifo_store[107][11] ),
    .A1(_04665_),
    .S(_04849_),
    .X(_04862_));
 sky130_fd_sc_hd__clkbuf_1 _09310_ (.A(_04862_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(\fifo0.fifo_store[107][12] ),
    .A1(_04751_),
    .S(_04849_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_1 _09312_ (.A(_04863_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(\fifo0.fifo_store[107][13] ),
    .A1(_04706_),
    .S(_04849_),
    .X(_04864_));
 sky130_fd_sc_hd__clkbuf_1 _09314_ (.A(_04864_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(\fifo0.fifo_store[107][14] ),
    .A1(_04754_),
    .S(_04849_),
    .X(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _09316_ (.A(_04865_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(\fifo0.fifo_store[107][15] ),
    .A1(_04756_),
    .S(_04849_),
    .X(_04866_));
 sky130_fd_sc_hd__clkbuf_1 _09318_ (.A(_04866_),
    .X(_00790_));
 sky130_fd_sc_hd__nor2_8 _09319_ (.A(_03965_),
    .B(_04629_),
    .Y(_04867_));
 sky130_fd_sc_hd__buf_8 _09320_ (.A(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(\fifo0.fifo_store[45][0] ),
    .A1(_04729_),
    .S(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _09322_ (.A(_04869_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(\fifo0.fifo_store[45][1] ),
    .A1(_04733_),
    .S(_04868_),
    .X(_04870_));
 sky130_fd_sc_hd__clkbuf_1 _09324_ (.A(_04870_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(\fifo0.fifo_store[45][2] ),
    .A1(_04735_),
    .S(_04868_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _09326_ (.A(_04871_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(\fifo0.fifo_store[45][3] ),
    .A1(_04737_),
    .S(_04868_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _09328_ (.A(_04872_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(\fifo0.fifo_store[45][4] ),
    .A1(_04739_),
    .S(_04868_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _09330_ (.A(_04873_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(\fifo0.fifo_store[45][5] ),
    .A1(_04656_),
    .S(_04868_),
    .X(_04874_));
 sky130_fd_sc_hd__clkbuf_1 _09332_ (.A(_04874_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(\fifo0.fifo_store[45][6] ),
    .A1(_04742_),
    .S(_04868_),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_1 _09334_ (.A(_04875_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(\fifo0.fifo_store[45][7] ),
    .A1(_04659_),
    .S(_04868_),
    .X(_04876_));
 sky130_fd_sc_hd__clkbuf_1 _09336_ (.A(_04876_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(\fifo0.fifo_store[45][8] ),
    .A1(_04745_),
    .S(_04868_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _09338_ (.A(_04877_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(\fifo0.fifo_store[45][9] ),
    .A1(_04747_),
    .S(_04868_),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_1 _09340_ (.A(_04878_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(\fifo0.fifo_store[45][10] ),
    .A1(_04663_),
    .S(_04867_),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _09342_ (.A(_04879_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(\fifo0.fifo_store[45][11] ),
    .A1(_04665_),
    .S(_04867_),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _09344_ (.A(_04880_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(\fifo0.fifo_store[45][12] ),
    .A1(_04751_),
    .S(_04867_),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _09346_ (.A(_04881_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _09347_ (.A0(\fifo0.fifo_store[45][13] ),
    .A1(_04706_),
    .S(_04867_),
    .X(_04882_));
 sky130_fd_sc_hd__clkbuf_1 _09348_ (.A(_04882_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(\fifo0.fifo_store[45][14] ),
    .A1(_04754_),
    .S(_04867_),
    .X(_04883_));
 sky130_fd_sc_hd__clkbuf_1 _09350_ (.A(_04883_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(\fifo0.fifo_store[45][15] ),
    .A1(_04756_),
    .S(_04867_),
    .X(_04884_));
 sky130_fd_sc_hd__clkbuf_1 _09352_ (.A(_04884_),
    .X(_00806_));
 sky130_fd_sc_hd__buf_4 _09353_ (.A(_03820_),
    .X(_04885_));
 sky130_fd_sc_hd__or2_1 _09354_ (.A(_04201_),
    .B(_04376_),
    .X(_04886_));
 sky130_fd_sc_hd__buf_4 _09355_ (.A(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_6 _09356_ (.A(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[126][0] ),
    .S(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_1 _09358_ (.A(_04889_),
    .X(_00807_));
 sky130_fd_sc_hd__buf_4 _09359_ (.A(_03828_),
    .X(_04890_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[126][1] ),
    .S(_04888_),
    .X(_04891_));
 sky130_fd_sc_hd__clkbuf_1 _09361_ (.A(_04891_),
    .X(_00808_));
 sky130_fd_sc_hd__buf_6 _09362_ (.A(_03831_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[126][2] ),
    .S(_04888_),
    .X(_04893_));
 sky130_fd_sc_hd__clkbuf_1 _09364_ (.A(_04893_),
    .X(_00809_));
 sky130_fd_sc_hd__buf_4 _09365_ (.A(_03833_),
    .X(_04894_));
 sky130_fd_sc_hd__mux2_1 _09366_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[126][3] ),
    .S(_04888_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_1 _09367_ (.A(_04895_),
    .X(_00810_));
 sky130_fd_sc_hd__buf_4 _09368_ (.A(_03835_),
    .X(_04896_));
 sky130_fd_sc_hd__mux2_1 _09369_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[126][4] ),
    .S(_04888_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_1 _09370_ (.A(_04897_),
    .X(_00811_));
 sky130_fd_sc_hd__buf_6 _09371_ (.A(_03838_),
    .X(_04898_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[126][5] ),
    .S(_04888_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_1 _09373_ (.A(_04899_),
    .X(_00812_));
 sky130_fd_sc_hd__buf_4 _09374_ (.A(_03840_),
    .X(_04900_));
 sky130_fd_sc_hd__mux2_1 _09375_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[126][6] ),
    .S(_04888_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_1 _09376_ (.A(_04901_),
    .X(_00813_));
 sky130_fd_sc_hd__clkbuf_8 _09377_ (.A(_03843_),
    .X(_04902_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[126][7] ),
    .S(_04888_),
    .X(_04903_));
 sky130_fd_sc_hd__clkbuf_1 _09379_ (.A(_04903_),
    .X(_00814_));
 sky130_fd_sc_hd__buf_6 _09380_ (.A(_03845_),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[126][8] ),
    .S(_04888_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_1 _09382_ (.A(_04905_),
    .X(_00815_));
 sky130_fd_sc_hd__buf_4 _09383_ (.A(_03847_),
    .X(_04906_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[126][9] ),
    .S(_04888_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_1 _09385_ (.A(_04907_),
    .X(_00816_));
 sky130_fd_sc_hd__buf_4 _09386_ (.A(_03850_),
    .X(_04908_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[126][10] ),
    .S(_04887_),
    .X(_04909_));
 sky130_fd_sc_hd__clkbuf_1 _09388_ (.A(_04909_),
    .X(_00817_));
 sky130_fd_sc_hd__buf_6 _09389_ (.A(_03853_),
    .X(_04910_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[126][11] ),
    .S(_04887_),
    .X(_04911_));
 sky130_fd_sc_hd__clkbuf_1 _09391_ (.A(_04911_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_6 _09392_ (.A(_03855_),
    .X(_04912_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[126][12] ),
    .S(_04887_),
    .X(_04913_));
 sky130_fd_sc_hd__clkbuf_1 _09394_ (.A(_04913_),
    .X(_00819_));
 sky130_fd_sc_hd__buf_6 _09395_ (.A(_03857_),
    .X(_04914_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[126][13] ),
    .S(_04887_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_1 _09397_ (.A(_04915_),
    .X(_00820_));
 sky130_fd_sc_hd__buf_6 _09398_ (.A(_03859_),
    .X(_04916_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[126][14] ),
    .S(_04887_),
    .X(_04917_));
 sky130_fd_sc_hd__clkbuf_1 _09400_ (.A(_04917_),
    .X(_00821_));
 sky130_fd_sc_hd__clkbuf_8 _09401_ (.A(_03861_),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[126][15] ),
    .S(_04887_),
    .X(_04919_));
 sky130_fd_sc_hd__clkbuf_1 _09403_ (.A(_04919_),
    .X(_00822_));
 sky130_fd_sc_hd__nor2_4 _09404_ (.A(_03965_),
    .B(_04376_),
    .Y(_04920_));
 sky130_fd_sc_hd__buf_6 _09405_ (.A(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(\fifo0.fifo_store[125][0] ),
    .A1(_04729_),
    .S(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__clkbuf_1 _09407_ (.A(_04922_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _09408_ (.A0(\fifo0.fifo_store[125][1] ),
    .A1(_04733_),
    .S(_04921_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_1 _09409_ (.A(_04923_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _09410_ (.A0(\fifo0.fifo_store[125][2] ),
    .A1(_04735_),
    .S(_04921_),
    .X(_04924_));
 sky130_fd_sc_hd__clkbuf_1 _09411_ (.A(_04924_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _09412_ (.A0(\fifo0.fifo_store[125][3] ),
    .A1(_04737_),
    .S(_04921_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_1 _09413_ (.A(_04925_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(\fifo0.fifo_store[125][4] ),
    .A1(_04739_),
    .S(_04921_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _09415_ (.A(_04926_),
    .X(_00827_));
 sky130_fd_sc_hd__buf_4 _09416_ (.A(_03838_),
    .X(_04927_));
 sky130_fd_sc_hd__mux2_1 _09417_ (.A0(\fifo0.fifo_store[125][5] ),
    .A1(_04927_),
    .S(_04921_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _09418_ (.A(_04928_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _09419_ (.A0(\fifo0.fifo_store[125][6] ),
    .A1(_04742_),
    .S(_04921_),
    .X(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _09420_ (.A(_04929_),
    .X(_00829_));
 sky130_fd_sc_hd__buf_4 _09421_ (.A(_03843_),
    .X(_04930_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(\fifo0.fifo_store[125][7] ),
    .A1(_04930_),
    .S(_04921_),
    .X(_04931_));
 sky130_fd_sc_hd__clkbuf_1 _09423_ (.A(_04931_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _09424_ (.A0(\fifo0.fifo_store[125][8] ),
    .A1(_04745_),
    .S(_04921_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _09425_ (.A(_04932_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _09426_ (.A0(\fifo0.fifo_store[125][9] ),
    .A1(_04747_),
    .S(_04921_),
    .X(_04933_));
 sky130_fd_sc_hd__clkbuf_1 _09427_ (.A(_04933_),
    .X(_00832_));
 sky130_fd_sc_hd__buf_4 _09428_ (.A(_03850_),
    .X(_04934_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(\fifo0.fifo_store[125][10] ),
    .A1(_04934_),
    .S(_04920_),
    .X(_04935_));
 sky130_fd_sc_hd__clkbuf_1 _09430_ (.A(_04935_),
    .X(_00833_));
 sky130_fd_sc_hd__buf_4 _09431_ (.A(_03853_),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _09432_ (.A0(\fifo0.fifo_store[125][11] ),
    .A1(_04936_),
    .S(_04920_),
    .X(_04937_));
 sky130_fd_sc_hd__clkbuf_1 _09433_ (.A(_04937_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _09434_ (.A0(\fifo0.fifo_store[125][12] ),
    .A1(_04751_),
    .S(_04920_),
    .X(_04938_));
 sky130_fd_sc_hd__clkbuf_1 _09435_ (.A(_04938_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _09436_ (.A0(\fifo0.fifo_store[125][13] ),
    .A1(_04706_),
    .S(_04920_),
    .X(_04939_));
 sky130_fd_sc_hd__clkbuf_1 _09437_ (.A(_04939_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(\fifo0.fifo_store[125][14] ),
    .A1(_04754_),
    .S(_04920_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_1 _09439_ (.A(_04940_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(\fifo0.fifo_store[125][15] ),
    .A1(_04756_),
    .S(_04920_),
    .X(_04941_));
 sky130_fd_sc_hd__clkbuf_1 _09441_ (.A(_04941_),
    .X(_00838_));
 sky130_fd_sc_hd__nor2_4 _09442_ (.A(_04032_),
    .B(_04145_),
    .Y(_04942_));
 sky130_fd_sc_hd__buf_6 _09443_ (.A(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(\fifo0.fifo_store[65][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_1 _09445_ (.A(_04944_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(\fifo0.fifo_store[65][1] ),
    .A1(_04733_),
    .S(_04943_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_1 _09447_ (.A(_04945_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _09448_ (.A0(\fifo0.fifo_store[65][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_04943_),
    .X(_04946_));
 sky130_fd_sc_hd__clkbuf_1 _09449_ (.A(_04946_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _09450_ (.A0(\fifo0.fifo_store[65][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_04943_),
    .X(_04947_));
 sky130_fd_sc_hd__clkbuf_1 _09451_ (.A(_04947_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(\fifo0.fifo_store[65][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_04943_),
    .X(_04948_));
 sky130_fd_sc_hd__clkbuf_1 _09453_ (.A(_04948_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(\fifo0.fifo_store[65][5] ),
    .A1(_04927_),
    .S(_04943_),
    .X(_04949_));
 sky130_fd_sc_hd__clkbuf_1 _09455_ (.A(_04949_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _09456_ (.A0(\fifo0.fifo_store[65][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_04943_),
    .X(_04950_));
 sky130_fd_sc_hd__clkbuf_1 _09457_ (.A(_04950_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(\fifo0.fifo_store[65][7] ),
    .A1(_04930_),
    .S(_04943_),
    .X(_04951_));
 sky130_fd_sc_hd__clkbuf_1 _09459_ (.A(_04951_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(\fifo0.fifo_store[65][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_04943_),
    .X(_04952_));
 sky130_fd_sc_hd__clkbuf_1 _09461_ (.A(_04952_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(\fifo0.fifo_store[65][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_04943_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _09463_ (.A(_04953_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(\fifo0.fifo_store[65][10] ),
    .A1(_04934_),
    .S(_04942_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_1 _09465_ (.A(_04954_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(\fifo0.fifo_store[65][11] ),
    .A1(_04936_),
    .S(_04942_),
    .X(_04955_));
 sky130_fd_sc_hd__clkbuf_1 _09467_ (.A(_04955_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _09468_ (.A0(\fifo0.fifo_store[65][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_04942_),
    .X(_04956_));
 sky130_fd_sc_hd__clkbuf_1 _09469_ (.A(_04956_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _09470_ (.A0(\fifo0.fifo_store[65][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_04942_),
    .X(_04957_));
 sky130_fd_sc_hd__clkbuf_1 _09471_ (.A(_04957_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _09472_ (.A0(\fifo0.fifo_store[65][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_04942_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_1 _09473_ (.A(_04958_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _09474_ (.A0(\fifo0.fifo_store[65][15] ),
    .A1(_04756_),
    .S(_04942_),
    .X(_04959_));
 sky130_fd_sc_hd__clkbuf_1 _09475_ (.A(_04959_),
    .X(_00854_));
 sky130_fd_sc_hd__nor2_4 _09476_ (.A(_03816_),
    .B(_04145_),
    .Y(_04960_));
 sky130_fd_sc_hd__buf_6 _09477_ (.A(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__mux2_1 _09478_ (.A0(\fifo0.fifo_store[64][0] ),
    .A1(_04729_),
    .S(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_1 _09479_ (.A(_04962_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(\fifo0.fifo_store[64][1] ),
    .A1(_04733_),
    .S(_04961_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_1 _09481_ (.A(_04963_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _09482_ (.A0(\fifo0.fifo_store[64][2] ),
    .A1(_04735_),
    .S(_04961_),
    .X(_04964_));
 sky130_fd_sc_hd__clkbuf_1 _09483_ (.A(_04964_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(\fifo0.fifo_store[64][3] ),
    .A1(_04737_),
    .S(_04961_),
    .X(_04965_));
 sky130_fd_sc_hd__clkbuf_1 _09485_ (.A(_04965_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _09486_ (.A0(\fifo0.fifo_store[64][4] ),
    .A1(_04739_),
    .S(_04961_),
    .X(_04966_));
 sky130_fd_sc_hd__clkbuf_1 _09487_ (.A(_04966_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _09488_ (.A0(\fifo0.fifo_store[64][5] ),
    .A1(_04927_),
    .S(_04961_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_1 _09489_ (.A(_04967_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _09490_ (.A0(\fifo0.fifo_store[64][6] ),
    .A1(_04742_),
    .S(_04961_),
    .X(_04968_));
 sky130_fd_sc_hd__clkbuf_1 _09491_ (.A(_04968_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(\fifo0.fifo_store[64][7] ),
    .A1(_04930_),
    .S(_04961_),
    .X(_04969_));
 sky130_fd_sc_hd__clkbuf_1 _09493_ (.A(_04969_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(\fifo0.fifo_store[64][8] ),
    .A1(_04745_),
    .S(_04961_),
    .X(_04970_));
 sky130_fd_sc_hd__clkbuf_1 _09495_ (.A(_04970_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _09496_ (.A0(\fifo0.fifo_store[64][9] ),
    .A1(_04747_),
    .S(_04961_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_1 _09497_ (.A(_04971_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(\fifo0.fifo_store[64][10] ),
    .A1(_04934_),
    .S(_04960_),
    .X(_04972_));
 sky130_fd_sc_hd__clkbuf_1 _09499_ (.A(_04972_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(\fifo0.fifo_store[64][11] ),
    .A1(_04936_),
    .S(_04960_),
    .X(_04973_));
 sky130_fd_sc_hd__clkbuf_1 _09501_ (.A(_04973_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _09502_ (.A0(\fifo0.fifo_store[64][12] ),
    .A1(_04751_),
    .S(_04960_),
    .X(_04974_));
 sky130_fd_sc_hd__clkbuf_1 _09503_ (.A(_04974_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(\fifo0.fifo_store[64][13] ),
    .A1(_04706_),
    .S(_04960_),
    .X(_04975_));
 sky130_fd_sc_hd__clkbuf_1 _09505_ (.A(_04975_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(\fifo0.fifo_store[64][14] ),
    .A1(_04754_),
    .S(_04960_),
    .X(_04976_));
 sky130_fd_sc_hd__clkbuf_1 _09507_ (.A(_04976_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _09508_ (.A0(\fifo0.fifo_store[64][15] ),
    .A1(_04756_),
    .S(_04960_),
    .X(_04977_));
 sky130_fd_sc_hd__clkbuf_1 _09509_ (.A(_04977_),
    .X(_00870_));
 sky130_fd_sc_hd__nor2_8 _09510_ (.A(_03990_),
    .B(_04172_),
    .Y(_04978_));
 sky130_fd_sc_hd__buf_12 _09511_ (.A(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(\fifo0.fifo_store[90][0] ),
    .A1(_04729_),
    .S(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__clkbuf_1 _09513_ (.A(_04980_),
    .X(_00871_));
 sky130_fd_sc_hd__buf_4 _09514_ (.A(_03872_),
    .X(_04981_));
 sky130_fd_sc_hd__mux2_1 _09515_ (.A0(\fifo0.fifo_store[90][1] ),
    .A1(_04981_),
    .S(_04979_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_1 _09516_ (.A(_04982_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _09517_ (.A0(\fifo0.fifo_store[90][2] ),
    .A1(_04735_),
    .S(_04979_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_1 _09518_ (.A(_04983_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _09519_ (.A0(\fifo0.fifo_store[90][3] ),
    .A1(_04737_),
    .S(_04979_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_1 _09520_ (.A(_04984_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(\fifo0.fifo_store[90][4] ),
    .A1(_04739_),
    .S(_04979_),
    .X(_04985_));
 sky130_fd_sc_hd__clkbuf_1 _09522_ (.A(_04985_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _09523_ (.A0(\fifo0.fifo_store[90][5] ),
    .A1(_04927_),
    .S(_04979_),
    .X(_04986_));
 sky130_fd_sc_hd__clkbuf_1 _09524_ (.A(_04986_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(\fifo0.fifo_store[90][6] ),
    .A1(_04742_),
    .S(_04979_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_1 _09526_ (.A(_04987_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _09527_ (.A0(\fifo0.fifo_store[90][7] ),
    .A1(_04930_),
    .S(_04979_),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_1 _09528_ (.A(_04988_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(\fifo0.fifo_store[90][8] ),
    .A1(_04745_),
    .S(_04979_),
    .X(_04989_));
 sky130_fd_sc_hd__clkbuf_1 _09530_ (.A(_04989_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(\fifo0.fifo_store[90][9] ),
    .A1(_04747_),
    .S(_04979_),
    .X(_04990_));
 sky130_fd_sc_hd__clkbuf_1 _09532_ (.A(_04990_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _09533_ (.A0(\fifo0.fifo_store[90][10] ),
    .A1(_04934_),
    .S(_04978_),
    .X(_04991_));
 sky130_fd_sc_hd__clkbuf_1 _09534_ (.A(_04991_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(\fifo0.fifo_store[90][11] ),
    .A1(_04936_),
    .S(_04978_),
    .X(_04992_));
 sky130_fd_sc_hd__clkbuf_1 _09536_ (.A(_04992_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(\fifo0.fifo_store[90][12] ),
    .A1(_04751_),
    .S(_04978_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_1 _09538_ (.A(_04993_),
    .X(_00883_));
 sky130_fd_sc_hd__clkbuf_4 _09539_ (.A(_03908_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _09540_ (.A0(\fifo0.fifo_store[90][13] ),
    .A1(_04994_),
    .S(_04978_),
    .X(_04995_));
 sky130_fd_sc_hd__clkbuf_1 _09541_ (.A(_04995_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _09542_ (.A0(\fifo0.fifo_store[90][14] ),
    .A1(_04754_),
    .S(_04978_),
    .X(_04996_));
 sky130_fd_sc_hd__clkbuf_1 _09543_ (.A(_04996_),
    .X(_00885_));
 sky130_fd_sc_hd__clkbuf_4 _09544_ (.A(_03914_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(\fifo0.fifo_store[90][15] ),
    .A1(_04997_),
    .S(_04978_),
    .X(_04998_));
 sky130_fd_sc_hd__clkbuf_1 _09546_ (.A(_04998_),
    .X(_00886_));
 sky130_fd_sc_hd__clkbuf_4 _09547_ (.A(_03821_),
    .X(_04999_));
 sky130_fd_sc_hd__or2_1 _09548_ (.A(_04170_),
    .B(_04627_),
    .X(_05000_));
 sky130_fd_sc_hd__buf_12 _09549_ (.A(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__nor2_8 _09550_ (.A(_03920_),
    .B(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__buf_12 _09551_ (.A(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(\fifo0.fifo_store[63][0] ),
    .A1(_04999_),
    .S(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__clkbuf_1 _09553_ (.A(_05004_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _09554_ (.A0(\fifo0.fifo_store[63][1] ),
    .A1(_04981_),
    .S(_05003_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_1 _09555_ (.A(_05005_),
    .X(_00888_));
 sky130_fd_sc_hd__clkbuf_8 _09556_ (.A(_03875_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(\fifo0.fifo_store[63][2] ),
    .A1(_05006_),
    .S(_05003_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _09558_ (.A(_05007_),
    .X(_00889_));
 sky130_fd_sc_hd__buf_4 _09559_ (.A(_03878_),
    .X(_05008_));
 sky130_fd_sc_hd__mux2_1 _09560_ (.A0(\fifo0.fifo_store[63][3] ),
    .A1(_05008_),
    .S(_05003_),
    .X(_05009_));
 sky130_fd_sc_hd__clkbuf_1 _09561_ (.A(_05009_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_4 _09562_ (.A(_03881_),
    .X(_05010_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(\fifo0.fifo_store[63][4] ),
    .A1(_05010_),
    .S(_05003_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_1 _09564_ (.A(_05011_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(\fifo0.fifo_store[63][5] ),
    .A1(_04927_),
    .S(_05003_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _09566_ (.A(_05012_),
    .X(_00892_));
 sky130_fd_sc_hd__buf_4 _09567_ (.A(_03887_),
    .X(_05013_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(\fifo0.fifo_store[63][6] ),
    .A1(_05013_),
    .S(_05003_),
    .X(_05014_));
 sky130_fd_sc_hd__clkbuf_1 _09569_ (.A(_05014_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(\fifo0.fifo_store[63][7] ),
    .A1(_04930_),
    .S(_05003_),
    .X(_05015_));
 sky130_fd_sc_hd__clkbuf_1 _09571_ (.A(_05015_),
    .X(_00894_));
 sky130_fd_sc_hd__buf_4 _09572_ (.A(_03893_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(\fifo0.fifo_store[63][8] ),
    .A1(_05016_),
    .S(_05003_),
    .X(_05017_));
 sky130_fd_sc_hd__clkbuf_1 _09574_ (.A(_05017_),
    .X(_00895_));
 sky130_fd_sc_hd__clkbuf_4 _09575_ (.A(_03896_),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _09576_ (.A0(\fifo0.fifo_store[63][9] ),
    .A1(_05018_),
    .S(_05003_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_1 _09577_ (.A(_05019_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _09578_ (.A0(\fifo0.fifo_store[63][10] ),
    .A1(_04934_),
    .S(_05002_),
    .X(_05020_));
 sky130_fd_sc_hd__clkbuf_1 _09579_ (.A(_05020_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _09580_ (.A0(\fifo0.fifo_store[63][11] ),
    .A1(_04936_),
    .S(_05002_),
    .X(_05021_));
 sky130_fd_sc_hd__clkbuf_1 _09581_ (.A(_05021_),
    .X(_00898_));
 sky130_fd_sc_hd__clkbuf_4 _09582_ (.A(_03905_),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(\fifo0.fifo_store[63][12] ),
    .A1(_05022_),
    .S(_05002_),
    .X(_05023_));
 sky130_fd_sc_hd__clkbuf_1 _09584_ (.A(_05023_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(\fifo0.fifo_store[63][13] ),
    .A1(_04994_),
    .S(_05002_),
    .X(_05024_));
 sky130_fd_sc_hd__clkbuf_1 _09586_ (.A(_05024_),
    .X(_00900_));
 sky130_fd_sc_hd__clkbuf_4 _09587_ (.A(_03911_),
    .X(_05025_));
 sky130_fd_sc_hd__mux2_1 _09588_ (.A0(\fifo0.fifo_store[63][14] ),
    .A1(_05025_),
    .S(_05002_),
    .X(_05026_));
 sky130_fd_sc_hd__clkbuf_1 _09589_ (.A(_05026_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(\fifo0.fifo_store[63][15] ),
    .A1(_04997_),
    .S(_05002_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_1 _09591_ (.A(_05027_),
    .X(_00902_));
 sky130_fd_sc_hd__or2_1 _09592_ (.A(_04201_),
    .B(_05001_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_4 _09593_ (.A(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_12 _09594_ (.A(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _09595_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[62][0] ),
    .S(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _09596_ (.A(_05031_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[62][1] ),
    .S(_05030_),
    .X(_05032_));
 sky130_fd_sc_hd__clkbuf_1 _09598_ (.A(_05032_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[62][2] ),
    .S(_05030_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _09600_ (.A(_05033_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[62][3] ),
    .S(_05030_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _09602_ (.A(_05034_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _09603_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[62][4] ),
    .S(_05030_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_1 _09604_ (.A(_05035_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[62][5] ),
    .S(_05030_),
    .X(_05036_));
 sky130_fd_sc_hd__clkbuf_1 _09606_ (.A(_05036_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _09607_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[62][6] ),
    .S(_05030_),
    .X(_05037_));
 sky130_fd_sc_hd__clkbuf_1 _09608_ (.A(_05037_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[62][7] ),
    .S(_05030_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _09610_ (.A(_05038_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _09611_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[62][8] ),
    .S(_05030_),
    .X(_05039_));
 sky130_fd_sc_hd__clkbuf_1 _09612_ (.A(_05039_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[62][9] ),
    .S(_05030_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_1 _09614_ (.A(_05040_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[62][10] ),
    .S(_05029_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_1 _09616_ (.A(_05041_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _09617_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[62][11] ),
    .S(_05029_),
    .X(_05042_));
 sky130_fd_sc_hd__clkbuf_1 _09618_ (.A(_05042_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _09619_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[62][12] ),
    .S(_05029_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _09620_ (.A(_05043_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _09621_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[62][13] ),
    .S(_05029_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _09622_ (.A(_05044_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[62][14] ),
    .S(_05029_),
    .X(_05045_));
 sky130_fd_sc_hd__clkbuf_1 _09624_ (.A(_05045_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[62][15] ),
    .S(_05029_),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_1 _09626_ (.A(_05046_),
    .X(_00918_));
 sky130_fd_sc_hd__nor2_8 _09627_ (.A(_03816_),
    .B(_04356_),
    .Y(_05047_));
 sky130_fd_sc_hd__buf_12 _09628_ (.A(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(\fifo0.fifo_store[8][0] ),
    .A1(_04999_),
    .S(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_1 _09630_ (.A(_05049_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(\fifo0.fifo_store[8][1] ),
    .A1(_04981_),
    .S(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _09632_ (.A(_05050_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(\fifo0.fifo_store[8][2] ),
    .A1(_05006_),
    .S(_05048_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _09634_ (.A(_05051_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(\fifo0.fifo_store[8][3] ),
    .A1(_05008_),
    .S(_05048_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _09636_ (.A(_05052_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(\fifo0.fifo_store[8][4] ),
    .A1(_05010_),
    .S(_05048_),
    .X(_05053_));
 sky130_fd_sc_hd__clkbuf_1 _09638_ (.A(_05053_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(\fifo0.fifo_store[8][5] ),
    .A1(_04927_),
    .S(_05048_),
    .X(_05054_));
 sky130_fd_sc_hd__clkbuf_1 _09640_ (.A(_05054_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(\fifo0.fifo_store[8][6] ),
    .A1(_05013_),
    .S(_05048_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _09642_ (.A(_05055_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _09643_ (.A0(\fifo0.fifo_store[8][7] ),
    .A1(_04930_),
    .S(_05048_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_1 _09644_ (.A(_05056_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(\fifo0.fifo_store[8][8] ),
    .A1(_05016_),
    .S(_05048_),
    .X(_05057_));
 sky130_fd_sc_hd__clkbuf_1 _09646_ (.A(_05057_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(\fifo0.fifo_store[8][9] ),
    .A1(_05018_),
    .S(_05048_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_1 _09648_ (.A(_05058_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(\fifo0.fifo_store[8][10] ),
    .A1(_04934_),
    .S(_05047_),
    .X(_05059_));
 sky130_fd_sc_hd__clkbuf_1 _09650_ (.A(_05059_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(\fifo0.fifo_store[8][11] ),
    .A1(_04936_),
    .S(_05047_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_05060_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(\fifo0.fifo_store[8][12] ),
    .A1(_05022_),
    .S(_05047_),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _09654_ (.A(_05061_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(\fifo0.fifo_store[8][13] ),
    .A1(_04994_),
    .S(_05047_),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _09656_ (.A(_05062_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _09657_ (.A0(\fifo0.fifo_store[8][14] ),
    .A1(_05025_),
    .S(_05047_),
    .X(_05063_));
 sky130_fd_sc_hd__clkbuf_1 _09658_ (.A(_05063_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _09659_ (.A0(\fifo0.fifo_store[8][15] ),
    .A1(_04997_),
    .S(_05047_),
    .X(_05064_));
 sky130_fd_sc_hd__clkbuf_1 _09660_ (.A(_05064_),
    .X(_00934_));
 sky130_fd_sc_hd__nor2_8 _09661_ (.A(_03965_),
    .B(_05001_),
    .Y(_05065_));
 sky130_fd_sc_hd__clkbuf_16 _09662_ (.A(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(\fifo0.fifo_store[61][0] ),
    .A1(_04999_),
    .S(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__clkbuf_1 _09664_ (.A(_05067_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(\fifo0.fifo_store[61][1] ),
    .A1(_04981_),
    .S(_05066_),
    .X(_05068_));
 sky130_fd_sc_hd__clkbuf_1 _09666_ (.A(_05068_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(\fifo0.fifo_store[61][2] ),
    .A1(_05006_),
    .S(_05066_),
    .X(_05069_));
 sky130_fd_sc_hd__clkbuf_1 _09668_ (.A(_05069_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(\fifo0.fifo_store[61][3] ),
    .A1(_05008_),
    .S(_05066_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _09670_ (.A(_05070_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(\fifo0.fifo_store[61][4] ),
    .A1(_05010_),
    .S(_05066_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_1 _09672_ (.A(_05071_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(\fifo0.fifo_store[61][5] ),
    .A1(_04927_),
    .S(_05066_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_1 _09674_ (.A(_05072_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(\fifo0.fifo_store[61][6] ),
    .A1(_05013_),
    .S(_05066_),
    .X(_05073_));
 sky130_fd_sc_hd__clkbuf_1 _09676_ (.A(_05073_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(\fifo0.fifo_store[61][7] ),
    .A1(_04930_),
    .S(_05066_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_1 _09678_ (.A(_05074_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(\fifo0.fifo_store[61][8] ),
    .A1(_05016_),
    .S(_05066_),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_1 _09680_ (.A(_05075_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(\fifo0.fifo_store[61][9] ),
    .A1(_05018_),
    .S(_05066_),
    .X(_05076_));
 sky130_fd_sc_hd__clkbuf_1 _09682_ (.A(_05076_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(\fifo0.fifo_store[61][10] ),
    .A1(_04934_),
    .S(_05065_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _09684_ (.A(_05077_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(\fifo0.fifo_store[61][11] ),
    .A1(_04936_),
    .S(_05065_),
    .X(_05078_));
 sky130_fd_sc_hd__clkbuf_1 _09686_ (.A(_05078_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(\fifo0.fifo_store[61][12] ),
    .A1(_05022_),
    .S(_05065_),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _09688_ (.A(_05079_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(\fifo0.fifo_store[61][13] ),
    .A1(_04994_),
    .S(_05065_),
    .X(_05080_));
 sky130_fd_sc_hd__clkbuf_1 _09690_ (.A(_05080_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(\fifo0.fifo_store[61][14] ),
    .A1(_05025_),
    .S(_05065_),
    .X(_05081_));
 sky130_fd_sc_hd__clkbuf_1 _09692_ (.A(_05081_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(\fifo0.fifo_store[61][15] ),
    .A1(_04997_),
    .S(_05065_),
    .X(_05082_));
 sky130_fd_sc_hd__clkbuf_1 _09694_ (.A(_05082_),
    .X(_00950_));
 sky130_fd_sc_hd__nor2_8 _09695_ (.A(_04277_),
    .B(_05001_),
    .Y(_05083_));
 sky130_fd_sc_hd__buf_12 _09696_ (.A(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__mux2_1 _09697_ (.A0(\fifo0.fifo_store[60][0] ),
    .A1(_04999_),
    .S(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__clkbuf_1 _09698_ (.A(_05085_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(\fifo0.fifo_store[60][1] ),
    .A1(_04981_),
    .S(_05084_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _09700_ (.A(_05086_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _09701_ (.A0(\fifo0.fifo_store[60][2] ),
    .A1(_05006_),
    .S(_05084_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_1 _09702_ (.A(_05087_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(\fifo0.fifo_store[60][3] ),
    .A1(_05008_),
    .S(_05084_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _09704_ (.A(_05088_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _09705_ (.A0(\fifo0.fifo_store[60][4] ),
    .A1(_05010_),
    .S(_05084_),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_1 _09706_ (.A(_05089_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _09707_ (.A0(\fifo0.fifo_store[60][5] ),
    .A1(_04927_),
    .S(_05084_),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _09708_ (.A(_05090_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _09709_ (.A0(\fifo0.fifo_store[60][6] ),
    .A1(_05013_),
    .S(_05084_),
    .X(_05091_));
 sky130_fd_sc_hd__clkbuf_1 _09710_ (.A(_05091_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(\fifo0.fifo_store[60][7] ),
    .A1(_04930_),
    .S(_05084_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _09712_ (.A(_05092_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(\fifo0.fifo_store[60][8] ),
    .A1(_05016_),
    .S(_05084_),
    .X(_05093_));
 sky130_fd_sc_hd__clkbuf_1 _09714_ (.A(_05093_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(\fifo0.fifo_store[60][9] ),
    .A1(_05018_),
    .S(_05084_),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _09716_ (.A(_05094_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(\fifo0.fifo_store[60][10] ),
    .A1(_04934_),
    .S(_05083_),
    .X(_05095_));
 sky130_fd_sc_hd__clkbuf_1 _09718_ (.A(_05095_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(\fifo0.fifo_store[60][11] ),
    .A1(_04936_),
    .S(_05083_),
    .X(_05096_));
 sky130_fd_sc_hd__clkbuf_1 _09720_ (.A(_05096_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(\fifo0.fifo_store[60][12] ),
    .A1(_05022_),
    .S(_05083_),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _09722_ (.A(_05097_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(\fifo0.fifo_store[60][13] ),
    .A1(_04994_),
    .S(_05083_),
    .X(_05098_));
 sky130_fd_sc_hd__clkbuf_1 _09724_ (.A(_05098_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(\fifo0.fifo_store[60][14] ),
    .A1(_05025_),
    .S(_05083_),
    .X(_05099_));
 sky130_fd_sc_hd__clkbuf_1 _09726_ (.A(_05099_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(\fifo0.fifo_store[60][15] ),
    .A1(_04997_),
    .S(_05083_),
    .X(_05100_));
 sky130_fd_sc_hd__clkbuf_1 _09728_ (.A(_05100_),
    .X(_00966_));
 sky130_fd_sc_hd__nor2_8 _09729_ (.A(_03815_),
    .B(_04172_),
    .Y(_05101_));
 sky130_fd_sc_hd__buf_12 _09730_ (.A(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _09731_ (.A0(\fifo0.fifo_store[88][0] ),
    .A1(_04999_),
    .S(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_1 _09732_ (.A(_05103_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(\fifo0.fifo_store[88][1] ),
    .A1(_04981_),
    .S(_05102_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _09734_ (.A(_05104_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(\fifo0.fifo_store[88][2] ),
    .A1(_05006_),
    .S(_05102_),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_1 _09736_ (.A(_05105_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(\fifo0.fifo_store[88][3] ),
    .A1(_05008_),
    .S(_05102_),
    .X(_05106_));
 sky130_fd_sc_hd__clkbuf_1 _09738_ (.A(_05106_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(\fifo0.fifo_store[88][4] ),
    .A1(_05010_),
    .S(_05102_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_1 _09740_ (.A(_05107_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(\fifo0.fifo_store[88][5] ),
    .A1(_04927_),
    .S(_05102_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _09742_ (.A(_05108_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(\fifo0.fifo_store[88][6] ),
    .A1(_05013_),
    .S(_05102_),
    .X(_05109_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_05109_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(\fifo0.fifo_store[88][7] ),
    .A1(_04930_),
    .S(_05102_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_1 _09746_ (.A(_05110_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\fifo0.fifo_store[88][8] ),
    .A1(_05016_),
    .S(_05102_),
    .X(_05111_));
 sky130_fd_sc_hd__clkbuf_1 _09748_ (.A(_05111_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(\fifo0.fifo_store[88][9] ),
    .A1(_05018_),
    .S(_05102_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(_05112_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _09751_ (.A0(\fifo0.fifo_store[88][10] ),
    .A1(_04934_),
    .S(_05101_),
    .X(_05113_));
 sky130_fd_sc_hd__clkbuf_1 _09752_ (.A(_05113_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _09753_ (.A0(\fifo0.fifo_store[88][11] ),
    .A1(_04936_),
    .S(_05101_),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_1 _09754_ (.A(_05114_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(\fifo0.fifo_store[88][12] ),
    .A1(_05022_),
    .S(_05101_),
    .X(_05115_));
 sky130_fd_sc_hd__clkbuf_1 _09756_ (.A(_05115_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _09757_ (.A0(\fifo0.fifo_store[88][13] ),
    .A1(_04994_),
    .S(_05101_),
    .X(_05116_));
 sky130_fd_sc_hd__clkbuf_1 _09758_ (.A(_05116_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _09759_ (.A0(\fifo0.fifo_store[88][14] ),
    .A1(_05025_),
    .S(_05101_),
    .X(_05117_));
 sky130_fd_sc_hd__clkbuf_1 _09760_ (.A(_05117_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(\fifo0.fifo_store[88][15] ),
    .A1(_04997_),
    .S(_05101_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_1 _09762_ (.A(_05118_),
    .X(_00982_));
 sky130_fd_sc_hd__nor2_4 _09763_ (.A(_03814_),
    .B(_03965_),
    .Y(_05119_));
 sky130_fd_sc_hd__buf_6 _09764_ (.A(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__mux2_1 _09765_ (.A0(\fifo0.fifo_store[5][0] ),
    .A1(_04999_),
    .S(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__clkbuf_1 _09766_ (.A(_05121_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(\fifo0.fifo_store[5][1] ),
    .A1(_04981_),
    .S(_05120_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _09768_ (.A(_05122_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(\fifo0.fifo_store[5][2] ),
    .A1(_05006_),
    .S(_05120_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _09770_ (.A(_05123_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(\fifo0.fifo_store[5][3] ),
    .A1(_05008_),
    .S(_05120_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_1 _09772_ (.A(_05124_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\fifo0.fifo_store[5][4] ),
    .A1(_05010_),
    .S(_05120_),
    .X(_05125_));
 sky130_fd_sc_hd__clkbuf_1 _09774_ (.A(_05125_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(\fifo0.fifo_store[5][5] ),
    .A1(_04927_),
    .S(_05120_),
    .X(_05126_));
 sky130_fd_sc_hd__clkbuf_1 _09776_ (.A(_05126_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _09777_ (.A0(\fifo0.fifo_store[5][6] ),
    .A1(_05013_),
    .S(_05120_),
    .X(_05127_));
 sky130_fd_sc_hd__clkbuf_1 _09778_ (.A(_05127_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(\fifo0.fifo_store[5][7] ),
    .A1(_04930_),
    .S(_05120_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _09780_ (.A(_05128_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(\fifo0.fifo_store[5][8] ),
    .A1(_05016_),
    .S(_05120_),
    .X(_05129_));
 sky130_fd_sc_hd__clkbuf_1 _09782_ (.A(_05129_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(\fifo0.fifo_store[5][9] ),
    .A1(_05018_),
    .S(_05120_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _09784_ (.A(_05130_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\fifo0.fifo_store[5][10] ),
    .A1(_04934_),
    .S(_05119_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_05131_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\fifo0.fifo_store[5][11] ),
    .A1(_04936_),
    .S(_05119_),
    .X(_05132_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_05132_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(\fifo0.fifo_store[5][12] ),
    .A1(_05022_),
    .S(_05119_),
    .X(_05133_));
 sky130_fd_sc_hd__clkbuf_1 _09790_ (.A(_05133_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(\fifo0.fifo_store[5][13] ),
    .A1(_04994_),
    .S(_05119_),
    .X(_05134_));
 sky130_fd_sc_hd__clkbuf_1 _09792_ (.A(_05134_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(\fifo0.fifo_store[5][14] ),
    .A1(_05025_),
    .S(_05119_),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_1 _09794_ (.A(_05135_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(\fifo0.fifo_store[5][15] ),
    .A1(_04997_),
    .S(_05119_),
    .X(_05136_));
 sky130_fd_sc_hd__clkbuf_1 _09796_ (.A(_05136_),
    .X(_00998_));
 sky130_fd_sc_hd__nor2_8 _09797_ (.A(_03990_),
    .B(_05001_),
    .Y(_05137_));
 sky130_fd_sc_hd__buf_8 _09798_ (.A(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_1 _09799_ (.A0(\fifo0.fifo_store[58][0] ),
    .A1(_04999_),
    .S(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_1 _09800_ (.A(_05139_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(\fifo0.fifo_store[58][1] ),
    .A1(_04981_),
    .S(_05138_),
    .X(_05140_));
 sky130_fd_sc_hd__clkbuf_1 _09802_ (.A(_05140_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(\fifo0.fifo_store[58][2] ),
    .A1(_05006_),
    .S(_05138_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _09804_ (.A(_05141_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(\fifo0.fifo_store[58][3] ),
    .A1(_05008_),
    .S(_05138_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _09806_ (.A(_05142_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _09807_ (.A0(\fifo0.fifo_store[58][4] ),
    .A1(_05010_),
    .S(_05138_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_1 _09808_ (.A(_05143_),
    .X(_01003_));
 sky130_fd_sc_hd__buf_4 _09809_ (.A(_03838_),
    .X(_05144_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(\fifo0.fifo_store[58][5] ),
    .A1(_05144_),
    .S(_05138_),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _09811_ (.A(_05145_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _09812_ (.A0(\fifo0.fifo_store[58][6] ),
    .A1(_05013_),
    .S(_05138_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_1 _09813_ (.A(_05146_),
    .X(_01005_));
 sky130_fd_sc_hd__clkbuf_4 _09814_ (.A(_03843_),
    .X(_05147_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(\fifo0.fifo_store[58][7] ),
    .A1(_05147_),
    .S(_05138_),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _09816_ (.A(_05148_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(\fifo0.fifo_store[58][8] ),
    .A1(_05016_),
    .S(_05138_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_1 _09818_ (.A(_05149_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(\fifo0.fifo_store[58][9] ),
    .A1(_05018_),
    .S(_05138_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _09820_ (.A(_05150_),
    .X(_01008_));
 sky130_fd_sc_hd__buf_2 _09821_ (.A(_03850_),
    .X(_05151_));
 sky130_fd_sc_hd__mux2_1 _09822_ (.A0(\fifo0.fifo_store[58][10] ),
    .A1(_05151_),
    .S(_05137_),
    .X(_05152_));
 sky130_fd_sc_hd__clkbuf_1 _09823_ (.A(_05152_),
    .X(_01009_));
 sky130_fd_sc_hd__buf_2 _09824_ (.A(_03853_),
    .X(_05153_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(\fifo0.fifo_store[58][11] ),
    .A1(_05153_),
    .S(_05137_),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_1 _09826_ (.A(_05154_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(\fifo0.fifo_store[58][12] ),
    .A1(_05022_),
    .S(_05137_),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_1 _09828_ (.A(_05155_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _09829_ (.A0(\fifo0.fifo_store[58][13] ),
    .A1(_04994_),
    .S(_05137_),
    .X(_05156_));
 sky130_fd_sc_hd__clkbuf_1 _09830_ (.A(_05156_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(\fifo0.fifo_store[58][14] ),
    .A1(_05025_),
    .S(_05137_),
    .X(_05157_));
 sky130_fd_sc_hd__clkbuf_1 _09832_ (.A(_05157_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(\fifo0.fifo_store[58][15] ),
    .A1(_04997_),
    .S(_05137_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_05158_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2_8 _09835_ (.A(_03868_),
    .B(_03920_),
    .Y(_05159_));
 sky130_fd_sc_hd__buf_12 _09836_ (.A(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(\fifo0.fifo_store[87][0] ),
    .A1(_04999_),
    .S(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__clkbuf_1 _09838_ (.A(_05161_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _09839_ (.A0(\fifo0.fifo_store[87][1] ),
    .A1(_04981_),
    .S(_05160_),
    .X(_05162_));
 sky130_fd_sc_hd__clkbuf_1 _09840_ (.A(_05162_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(\fifo0.fifo_store[87][2] ),
    .A1(_05006_),
    .S(_05160_),
    .X(_05163_));
 sky130_fd_sc_hd__clkbuf_1 _09842_ (.A(_05163_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(\fifo0.fifo_store[87][3] ),
    .A1(_05008_),
    .S(_05160_),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_1 _09844_ (.A(_05164_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(\fifo0.fifo_store[87][4] ),
    .A1(_05010_),
    .S(_05160_),
    .X(_05165_));
 sky130_fd_sc_hd__clkbuf_1 _09846_ (.A(_05165_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(\fifo0.fifo_store[87][5] ),
    .A1(_05144_),
    .S(_05160_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _09848_ (.A(_05166_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(\fifo0.fifo_store[87][6] ),
    .A1(_05013_),
    .S(_05160_),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _09850_ (.A(_05167_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(\fifo0.fifo_store[87][7] ),
    .A1(_05147_),
    .S(_05160_),
    .X(_05168_));
 sky130_fd_sc_hd__clkbuf_1 _09852_ (.A(_05168_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(\fifo0.fifo_store[87][8] ),
    .A1(_05016_),
    .S(_05160_),
    .X(_05169_));
 sky130_fd_sc_hd__clkbuf_1 _09854_ (.A(_05169_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _09855_ (.A0(\fifo0.fifo_store[87][9] ),
    .A1(_05018_),
    .S(_05160_),
    .X(_05170_));
 sky130_fd_sc_hd__clkbuf_1 _09856_ (.A(_05170_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _09857_ (.A0(\fifo0.fifo_store[87][10] ),
    .A1(_05151_),
    .S(_05159_),
    .X(_05171_));
 sky130_fd_sc_hd__clkbuf_1 _09858_ (.A(_05171_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _09859_ (.A0(\fifo0.fifo_store[87][11] ),
    .A1(_05153_),
    .S(_05159_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_1 _09860_ (.A(_05172_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _09861_ (.A0(\fifo0.fifo_store[87][12] ),
    .A1(_05022_),
    .S(_05159_),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_1 _09862_ (.A(_05173_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _09863_ (.A0(\fifo0.fifo_store[87][13] ),
    .A1(_04994_),
    .S(_05159_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_1 _09864_ (.A(_05174_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _09865_ (.A0(\fifo0.fifo_store[87][14] ),
    .A1(_05025_),
    .S(_05159_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_1 _09866_ (.A(_05175_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(\fifo0.fifo_store[87][15] ),
    .A1(_04997_),
    .S(_05159_),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_1 _09868_ (.A(_05176_),
    .X(_01030_));
 sky130_fd_sc_hd__nor2_8 _09869_ (.A(_04032_),
    .B(_05001_),
    .Y(_05177_));
 sky130_fd_sc_hd__buf_8 _09870_ (.A(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__mux2_1 _09871_ (.A0(\fifo0.fifo_store[57][0] ),
    .A1(_04999_),
    .S(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_1 _09872_ (.A(_05179_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(\fifo0.fifo_store[57][1] ),
    .A1(_04981_),
    .S(_05178_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_1 _09874_ (.A(_05180_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _09875_ (.A0(\fifo0.fifo_store[57][2] ),
    .A1(_05006_),
    .S(_05178_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _09876_ (.A(_05181_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(\fifo0.fifo_store[57][3] ),
    .A1(_05008_),
    .S(_05178_),
    .X(_05182_));
 sky130_fd_sc_hd__clkbuf_1 _09878_ (.A(_05182_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(\fifo0.fifo_store[57][4] ),
    .A1(_05010_),
    .S(_05178_),
    .X(_05183_));
 sky130_fd_sc_hd__clkbuf_1 _09880_ (.A(_05183_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(\fifo0.fifo_store[57][5] ),
    .A1(_05144_),
    .S(_05178_),
    .X(_05184_));
 sky130_fd_sc_hd__clkbuf_1 _09882_ (.A(_05184_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(\fifo0.fifo_store[57][6] ),
    .A1(_05013_),
    .S(_05178_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_1 _09884_ (.A(_05185_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(\fifo0.fifo_store[57][7] ),
    .A1(_05147_),
    .S(_05178_),
    .X(_05186_));
 sky130_fd_sc_hd__clkbuf_1 _09886_ (.A(_05186_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _09887_ (.A0(\fifo0.fifo_store[57][8] ),
    .A1(_05016_),
    .S(_05178_),
    .X(_05187_));
 sky130_fd_sc_hd__clkbuf_1 _09888_ (.A(_05187_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _09889_ (.A0(\fifo0.fifo_store[57][9] ),
    .A1(_05018_),
    .S(_05178_),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_1 _09890_ (.A(_05188_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(\fifo0.fifo_store[57][10] ),
    .A1(_05151_),
    .S(_05177_),
    .X(_05189_));
 sky130_fd_sc_hd__clkbuf_1 _09892_ (.A(_05189_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _09893_ (.A0(\fifo0.fifo_store[57][11] ),
    .A1(_05153_),
    .S(_05177_),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_1 _09894_ (.A(_05190_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _09895_ (.A0(\fifo0.fifo_store[57][12] ),
    .A1(_05022_),
    .S(_05177_),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_1 _09896_ (.A(_05191_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _09897_ (.A0(\fifo0.fifo_store[57][13] ),
    .A1(_04994_),
    .S(_05177_),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _09898_ (.A(_05192_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _09899_ (.A0(\fifo0.fifo_store[57][14] ),
    .A1(_05025_),
    .S(_05177_),
    .X(_05193_));
 sky130_fd_sc_hd__clkbuf_1 _09900_ (.A(_05193_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _09901_ (.A0(\fifo0.fifo_store[57][15] ),
    .A1(_04997_),
    .S(_05177_),
    .X(_05194_));
 sky130_fd_sc_hd__clkbuf_1 _09902_ (.A(_05194_),
    .X(_01046_));
 sky130_fd_sc_hd__nor2_8 _09903_ (.A(_03815_),
    .B(_05001_),
    .Y(_05195_));
 sky130_fd_sc_hd__buf_8 _09904_ (.A(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _09905_ (.A0(\fifo0.fifo_store[56][0] ),
    .A1(_04999_),
    .S(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_1 _09906_ (.A(_05197_),
    .X(_01047_));
 sky130_fd_sc_hd__buf_4 _09907_ (.A(_03872_),
    .X(_05198_));
 sky130_fd_sc_hd__mux2_1 _09908_ (.A0(\fifo0.fifo_store[56][1] ),
    .A1(_05198_),
    .S(_05196_),
    .X(_05199_));
 sky130_fd_sc_hd__clkbuf_1 _09909_ (.A(_05199_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _09910_ (.A0(\fifo0.fifo_store[56][2] ),
    .A1(_05006_),
    .S(_05196_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_1 _09911_ (.A(_05200_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(\fifo0.fifo_store[56][3] ),
    .A1(_05008_),
    .S(_05196_),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_1 _09913_ (.A(_05201_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _09914_ (.A0(\fifo0.fifo_store[56][4] ),
    .A1(_05010_),
    .S(_05196_),
    .X(_05202_));
 sky130_fd_sc_hd__clkbuf_1 _09915_ (.A(_05202_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(\fifo0.fifo_store[56][5] ),
    .A1(_05144_),
    .S(_05196_),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_1 _09917_ (.A(_05203_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(\fifo0.fifo_store[56][6] ),
    .A1(_05013_),
    .S(_05196_),
    .X(_05204_));
 sky130_fd_sc_hd__clkbuf_1 _09919_ (.A(_05204_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(\fifo0.fifo_store[56][7] ),
    .A1(_05147_),
    .S(_05196_),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_1 _09921_ (.A(_05205_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(\fifo0.fifo_store[56][8] ),
    .A1(_05016_),
    .S(_05196_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _09923_ (.A(_05206_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(\fifo0.fifo_store[56][9] ),
    .A1(_05018_),
    .S(_05196_),
    .X(_05207_));
 sky130_fd_sc_hd__clkbuf_1 _09925_ (.A(_05207_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _09926_ (.A0(\fifo0.fifo_store[56][10] ),
    .A1(_05151_),
    .S(_05195_),
    .X(_05208_));
 sky130_fd_sc_hd__clkbuf_1 _09927_ (.A(_05208_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(\fifo0.fifo_store[56][11] ),
    .A1(_05153_),
    .S(_05195_),
    .X(_05209_));
 sky130_fd_sc_hd__clkbuf_1 _09929_ (.A(_05209_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _09930_ (.A0(\fifo0.fifo_store[56][12] ),
    .A1(_05022_),
    .S(_05195_),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_1 _09931_ (.A(_05210_),
    .X(_01059_));
 sky130_fd_sc_hd__clkbuf_4 _09932_ (.A(_03908_),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(\fifo0.fifo_store[56][13] ),
    .A1(_05211_),
    .S(_05195_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_1 _09934_ (.A(_05212_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(\fifo0.fifo_store[56][14] ),
    .A1(_05025_),
    .S(_05195_),
    .X(_05213_));
 sky130_fd_sc_hd__clkbuf_1 _09936_ (.A(_05213_),
    .X(_01061_));
 sky130_fd_sc_hd__clkbuf_4 _09937_ (.A(_03914_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(\fifo0.fifo_store[56][15] ),
    .A1(_05214_),
    .S(_05195_),
    .X(_05215_));
 sky130_fd_sc_hd__clkbuf_1 _09939_ (.A(_05215_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _09940_ (.A(_03868_),
    .B(_03943_),
    .X(_05216_));
 sky130_fd_sc_hd__buf_4 _09941_ (.A(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__buf_12 _09942_ (.A(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__mux2_1 _09943_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[86][0] ),
    .S(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__clkbuf_1 _09944_ (.A(_05219_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _09945_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[86][1] ),
    .S(_05218_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_1 _09946_ (.A(_05220_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[86][2] ),
    .S(_05218_),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_1 _09948_ (.A(_05221_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[86][3] ),
    .S(_05218_),
    .X(_05222_));
 sky130_fd_sc_hd__clkbuf_1 _09950_ (.A(_05222_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[86][4] ),
    .S(_05218_),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_1 _09952_ (.A(_05223_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[86][5] ),
    .S(_05218_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_05224_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[86][6] ),
    .S(_05218_),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _09956_ (.A(_05225_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[86][7] ),
    .S(_05218_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _09958_ (.A(_05226_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[86][8] ),
    .S(_05218_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _09960_ (.A(_05227_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[86][9] ),
    .S(_05218_),
    .X(_05228_));
 sky130_fd_sc_hd__clkbuf_1 _09962_ (.A(_05228_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[86][10] ),
    .S(_05217_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _09964_ (.A(_05229_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[86][11] ),
    .S(_05217_),
    .X(_05230_));
 sky130_fd_sc_hd__clkbuf_1 _09966_ (.A(_05230_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[86][12] ),
    .S(_05217_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _09968_ (.A(_05231_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[86][13] ),
    .S(_05217_),
    .X(_05232_));
 sky130_fd_sc_hd__clkbuf_1 _09970_ (.A(_05232_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[86][14] ),
    .S(_05217_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _09972_ (.A(_05233_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[86][15] ),
    .S(_05217_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_1 _09974_ (.A(_05234_),
    .X(_01078_));
 sky130_fd_sc_hd__clkbuf_4 _09975_ (.A(_03821_),
    .X(_05235_));
 sky130_fd_sc_hd__nor2_8 _09976_ (.A(_03920_),
    .B(_04690_),
    .Y(_05236_));
 sky130_fd_sc_hd__buf_12 _09977_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(\fifo0.fifo_store[55][0] ),
    .A1(_05235_),
    .S(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__clkbuf_1 _09979_ (.A(_05238_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _09980_ (.A0(\fifo0.fifo_store[55][1] ),
    .A1(_05198_),
    .S(_05237_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_1 _09981_ (.A(_05239_),
    .X(_01080_));
 sky130_fd_sc_hd__buf_4 _09982_ (.A(_03875_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_1 _09983_ (.A0(\fifo0.fifo_store[55][2] ),
    .A1(_05240_),
    .S(_05237_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _09984_ (.A(_05241_),
    .X(_01081_));
 sky130_fd_sc_hd__clkbuf_4 _09985_ (.A(_03878_),
    .X(_05242_));
 sky130_fd_sc_hd__mux2_1 _09986_ (.A0(\fifo0.fifo_store[55][3] ),
    .A1(_05242_),
    .S(_05237_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _09987_ (.A(_05243_),
    .X(_01082_));
 sky130_fd_sc_hd__clkbuf_4 _09988_ (.A(_03881_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_1 _09989_ (.A0(\fifo0.fifo_store[55][4] ),
    .A1(_05244_),
    .S(_05237_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_1 _09990_ (.A(_05245_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(\fifo0.fifo_store[55][5] ),
    .A1(_05144_),
    .S(_05237_),
    .X(_05246_));
 sky130_fd_sc_hd__clkbuf_1 _09992_ (.A(_05246_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _09993_ (.A(_03887_),
    .X(_05247_));
 sky130_fd_sc_hd__mux2_1 _09994_ (.A0(\fifo0.fifo_store[55][6] ),
    .A1(_05247_),
    .S(_05237_),
    .X(_05248_));
 sky130_fd_sc_hd__clkbuf_1 _09995_ (.A(_05248_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(\fifo0.fifo_store[55][7] ),
    .A1(_05147_),
    .S(_05237_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _09997_ (.A(_05249_),
    .X(_01086_));
 sky130_fd_sc_hd__clkbuf_4 _09998_ (.A(_03893_),
    .X(_05250_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(\fifo0.fifo_store[55][8] ),
    .A1(_05250_),
    .S(_05237_),
    .X(_05251_));
 sky130_fd_sc_hd__clkbuf_1 _10000_ (.A(_05251_),
    .X(_01087_));
 sky130_fd_sc_hd__clkbuf_4 _10001_ (.A(_03896_),
    .X(_05252_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(\fifo0.fifo_store[55][9] ),
    .A1(_05252_),
    .S(_05237_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _10003_ (.A(_05253_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(\fifo0.fifo_store[55][10] ),
    .A1(_05151_),
    .S(_05236_),
    .X(_05254_));
 sky130_fd_sc_hd__clkbuf_1 _10005_ (.A(_05254_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(\fifo0.fifo_store[55][11] ),
    .A1(_05153_),
    .S(_05236_),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_1 _10007_ (.A(_05255_),
    .X(_01090_));
 sky130_fd_sc_hd__buf_4 _10008_ (.A(_03905_),
    .X(_05256_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(\fifo0.fifo_store[55][12] ),
    .A1(_05256_),
    .S(_05236_),
    .X(_05257_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_05257_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(\fifo0.fifo_store[55][13] ),
    .A1(_05211_),
    .S(_05236_),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_1 _10012_ (.A(_05258_),
    .X(_01092_));
 sky130_fd_sc_hd__buf_4 _10013_ (.A(_03911_),
    .X(_05259_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(\fifo0.fifo_store[55][14] ),
    .A1(_05259_),
    .S(_05236_),
    .X(_05260_));
 sky130_fd_sc_hd__clkbuf_1 _10015_ (.A(_05260_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(\fifo0.fifo_store[55][15] ),
    .A1(_05214_),
    .S(_05236_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _10017_ (.A(_05261_),
    .X(_01094_));
 sky130_fd_sc_hd__nor2_8 _10018_ (.A(_03868_),
    .B(_03965_),
    .Y(_05262_));
 sky130_fd_sc_hd__buf_12 _10019_ (.A(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(\fifo0.fifo_store[85][0] ),
    .A1(_05235_),
    .S(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _10021_ (.A(_05264_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(\fifo0.fifo_store[85][1] ),
    .A1(_05198_),
    .S(_05263_),
    .X(_05265_));
 sky130_fd_sc_hd__clkbuf_1 _10023_ (.A(_05265_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(\fifo0.fifo_store[85][2] ),
    .A1(_05240_),
    .S(_05263_),
    .X(_05266_));
 sky130_fd_sc_hd__clkbuf_1 _10025_ (.A(_05266_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(\fifo0.fifo_store[85][3] ),
    .A1(_05242_),
    .S(_05263_),
    .X(_05267_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_05267_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(\fifo0.fifo_store[85][4] ),
    .A1(_05244_),
    .S(_05263_),
    .X(_05268_));
 sky130_fd_sc_hd__clkbuf_1 _10029_ (.A(_05268_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(\fifo0.fifo_store[85][5] ),
    .A1(_05144_),
    .S(_05263_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_1 _10031_ (.A(_05269_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(\fifo0.fifo_store[85][6] ),
    .A1(_05247_),
    .S(_05263_),
    .X(_05270_));
 sky130_fd_sc_hd__clkbuf_1 _10033_ (.A(_05270_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\fifo0.fifo_store[85][7] ),
    .A1(_05147_),
    .S(_05263_),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_1 _10035_ (.A(_05271_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(\fifo0.fifo_store[85][8] ),
    .A1(_05250_),
    .S(_05263_),
    .X(_05272_));
 sky130_fd_sc_hd__clkbuf_1 _10037_ (.A(_05272_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\fifo0.fifo_store[85][9] ),
    .A1(_05252_),
    .S(_05263_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _10039_ (.A(_05273_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(\fifo0.fifo_store[85][10] ),
    .A1(_05151_),
    .S(_05262_),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_1 _10041_ (.A(_05274_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(\fifo0.fifo_store[85][11] ),
    .A1(_05153_),
    .S(_05262_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _10043_ (.A(_05275_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _10044_ (.A0(\fifo0.fifo_store[85][12] ),
    .A1(_05256_),
    .S(_05262_),
    .X(_05276_));
 sky130_fd_sc_hd__clkbuf_1 _10045_ (.A(_05276_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\fifo0.fifo_store[85][13] ),
    .A1(_05211_),
    .S(_05262_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_1 _10047_ (.A(_05277_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(\fifo0.fifo_store[85][14] ),
    .A1(_05259_),
    .S(_05262_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_1 _10049_ (.A(_05278_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(\fifo0.fifo_store[85][15] ),
    .A1(_05214_),
    .S(_05262_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_1 _10051_ (.A(_05279_),
    .X(_01110_));
 sky130_fd_sc_hd__or2_1 _10052_ (.A(_04201_),
    .B(_04690_),
    .X(_05280_));
 sky130_fd_sc_hd__buf_4 _10053_ (.A(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__buf_12 _10054_ (.A(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[54][0] ),
    .S(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _10056_ (.A(_05283_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[54][1] ),
    .S(_05282_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_05284_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[54][2] ),
    .S(_05282_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _10060_ (.A(_05285_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _10061_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[54][3] ),
    .S(_05282_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_1 _10062_ (.A(_05286_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[54][4] ),
    .S(_05282_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_1 _10064_ (.A(_05287_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _10065_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[54][5] ),
    .S(_05282_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _10066_ (.A(_05288_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _10067_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[54][6] ),
    .S(_05282_),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_1 _10068_ (.A(_05289_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[54][7] ),
    .S(_05282_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_1 _10070_ (.A(_05290_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[54][8] ),
    .S(_05282_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_1 _10072_ (.A(_05291_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[54][9] ),
    .S(_05282_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _10074_ (.A(_05292_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[54][10] ),
    .S(_05281_),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_05293_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[54][11] ),
    .S(_05281_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _10078_ (.A(_05294_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[54][12] ),
    .S(_05281_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_1 _10080_ (.A(_05295_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[54][13] ),
    .S(_05281_),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_1 _10082_ (.A(_05296_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[54][14] ),
    .S(_05281_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_1 _10084_ (.A(_05297_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[54][15] ),
    .S(_05281_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _10086_ (.A(_05298_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _10087_ (.A(_03868_),
    .B(_04010_),
    .X(_05299_));
 sky130_fd_sc_hd__buf_4 _10088_ (.A(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__buf_12 _10089_ (.A(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[84][0] ),
    .S(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_1 _10091_ (.A(_05302_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[84][1] ),
    .S(_05301_),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_1 _10093_ (.A(_05303_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[84][2] ),
    .S(_05301_),
    .X(_05304_));
 sky130_fd_sc_hd__clkbuf_1 _10095_ (.A(_05304_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _10096_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[84][3] ),
    .S(_05301_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _10097_ (.A(_05305_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _10098_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[84][4] ),
    .S(_05301_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _10099_ (.A(_05306_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[84][5] ),
    .S(_05301_),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_1 _10101_ (.A(_05307_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _10102_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[84][6] ),
    .S(_05301_),
    .X(_05308_));
 sky130_fd_sc_hd__clkbuf_1 _10103_ (.A(_05308_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _10104_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[84][7] ),
    .S(_05301_),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _10105_ (.A(_05309_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _10106_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[84][8] ),
    .S(_05301_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_1 _10107_ (.A(_05310_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _10108_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[84][9] ),
    .S(_05301_),
    .X(_05311_));
 sky130_fd_sc_hd__clkbuf_1 _10109_ (.A(_05311_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _10110_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[84][10] ),
    .S(_05300_),
    .X(_05312_));
 sky130_fd_sc_hd__clkbuf_1 _10111_ (.A(_05312_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[84][11] ),
    .S(_05300_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_1 _10113_ (.A(_05313_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[84][12] ),
    .S(_05300_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_1 _10115_ (.A(_05314_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[84][13] ),
    .S(_05300_),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_1 _10117_ (.A(_05315_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[84][14] ),
    .S(_05300_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _10119_ (.A(_05316_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[84][15] ),
    .S(_05300_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_1 _10121_ (.A(_05317_),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_8 _10122_ (.A(_03965_),
    .B(_04690_),
    .Y(_05318_));
 sky130_fd_sc_hd__buf_12 _10123_ (.A(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(\fifo0.fifo_store[53][0] ),
    .A1(_05235_),
    .S(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _10125_ (.A(_05320_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(\fifo0.fifo_store[53][1] ),
    .A1(_05198_),
    .S(_05319_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_1 _10127_ (.A(_05321_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(\fifo0.fifo_store[53][2] ),
    .A1(_05240_),
    .S(_05319_),
    .X(_05322_));
 sky130_fd_sc_hd__clkbuf_1 _10129_ (.A(_05322_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\fifo0.fifo_store[53][3] ),
    .A1(_05242_),
    .S(_05319_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_1 _10131_ (.A(_05323_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(\fifo0.fifo_store[53][4] ),
    .A1(_05244_),
    .S(_05319_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _10133_ (.A(_05324_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\fifo0.fifo_store[53][5] ),
    .A1(_05144_),
    .S(_05319_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _10135_ (.A(_05325_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\fifo0.fifo_store[53][6] ),
    .A1(_05247_),
    .S(_05319_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_1 _10137_ (.A(_05326_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\fifo0.fifo_store[53][7] ),
    .A1(_05147_),
    .S(_05319_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _10139_ (.A(_05327_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(\fifo0.fifo_store[53][8] ),
    .A1(_05250_),
    .S(_05319_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_1 _10141_ (.A(_05328_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(\fifo0.fifo_store[53][9] ),
    .A1(_05252_),
    .S(_05319_),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _10143_ (.A(_05329_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _10144_ (.A0(\fifo0.fifo_store[53][10] ),
    .A1(_05151_),
    .S(_05318_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _10145_ (.A(_05330_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(\fifo0.fifo_store[53][11] ),
    .A1(_05153_),
    .S(_05318_),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _10147_ (.A(_05331_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(\fifo0.fifo_store[53][12] ),
    .A1(_05256_),
    .S(_05318_),
    .X(_05332_));
 sky130_fd_sc_hd__clkbuf_1 _10149_ (.A(_05332_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\fifo0.fifo_store[53][13] ),
    .A1(_05211_),
    .S(_05318_),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _10151_ (.A(_05333_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(\fifo0.fifo_store[53][14] ),
    .A1(_05259_),
    .S(_05318_),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_1 _10153_ (.A(_05334_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(\fifo0.fifo_store[53][15] ),
    .A1(_05214_),
    .S(_05318_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _10155_ (.A(_05335_),
    .X(_01158_));
 sky130_fd_sc_hd__nor2_8 _10156_ (.A(_04277_),
    .B(_04690_),
    .Y(_05336_));
 sky130_fd_sc_hd__buf_12 _10157_ (.A(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _10158_ (.A0(\fifo0.fifo_store[52][0] ),
    .A1(_05235_),
    .S(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _10159_ (.A(_05338_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(\fifo0.fifo_store[52][1] ),
    .A1(_05198_),
    .S(_05337_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _10161_ (.A(_05339_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _10162_ (.A0(\fifo0.fifo_store[52][2] ),
    .A1(_05240_),
    .S(_05337_),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _10163_ (.A(_05340_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(\fifo0.fifo_store[52][3] ),
    .A1(_05242_),
    .S(_05337_),
    .X(_05341_));
 sky130_fd_sc_hd__clkbuf_1 _10165_ (.A(_05341_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(\fifo0.fifo_store[52][4] ),
    .A1(_05244_),
    .S(_05337_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_1 _10167_ (.A(_05342_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _10168_ (.A0(\fifo0.fifo_store[52][5] ),
    .A1(_05144_),
    .S(_05337_),
    .X(_05343_));
 sky130_fd_sc_hd__clkbuf_1 _10169_ (.A(_05343_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(\fifo0.fifo_store[52][6] ),
    .A1(_05247_),
    .S(_05337_),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_1 _10171_ (.A(_05344_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(\fifo0.fifo_store[52][7] ),
    .A1(_05147_),
    .S(_05337_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _10173_ (.A(_05345_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(\fifo0.fifo_store[52][8] ),
    .A1(_05250_),
    .S(_05337_),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_1 _10175_ (.A(_05346_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(\fifo0.fifo_store[52][9] ),
    .A1(_05252_),
    .S(_05337_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _10177_ (.A(_05347_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _10178_ (.A0(\fifo0.fifo_store[52][10] ),
    .A1(_05151_),
    .S(_05336_),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _10179_ (.A(_05348_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(\fifo0.fifo_store[52][11] ),
    .A1(_05153_),
    .S(_05336_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _10181_ (.A(_05349_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(\fifo0.fifo_store[52][12] ),
    .A1(_05256_),
    .S(_05336_),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_1 _10183_ (.A(_05350_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(\fifo0.fifo_store[52][13] ),
    .A1(_05211_),
    .S(_05336_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _10185_ (.A(_05351_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(\fifo0.fifo_store[52][14] ),
    .A1(_05259_),
    .S(_05336_),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _10187_ (.A(_05352_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(\fifo0.fifo_store[52][15] ),
    .A1(_05214_),
    .S(_05336_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _10189_ (.A(_05353_),
    .X(_01174_));
 sky130_fd_sc_hd__nor2_8 _10190_ (.A(_03868_),
    .B(_04053_),
    .Y(_05354_));
 sky130_fd_sc_hd__buf_6 _10191_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(\fifo0.fifo_store[83][0] ),
    .A1(_05235_),
    .S(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_05356_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(\fifo0.fifo_store[83][1] ),
    .A1(_05198_),
    .S(_05355_),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_05357_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(\fifo0.fifo_store[83][2] ),
    .A1(_05240_),
    .S(_05355_),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _10197_ (.A(_05358_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(\fifo0.fifo_store[83][3] ),
    .A1(_05242_),
    .S(_05355_),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _10199_ (.A(_05359_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(\fifo0.fifo_store[83][4] ),
    .A1(_05244_),
    .S(_05355_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_05360_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(\fifo0.fifo_store[83][5] ),
    .A1(_05144_),
    .S(_05355_),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _10203_ (.A(_05361_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(\fifo0.fifo_store[83][6] ),
    .A1(_05247_),
    .S(_05355_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _10205_ (.A(_05362_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\fifo0.fifo_store[83][7] ),
    .A1(_05147_),
    .S(_05355_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _10207_ (.A(_05363_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(\fifo0.fifo_store[83][8] ),
    .A1(_05250_),
    .S(_05355_),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(_05364_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(\fifo0.fifo_store[83][9] ),
    .A1(_05252_),
    .S(_05355_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _10211_ (.A(_05365_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(\fifo0.fifo_store[83][10] ),
    .A1(_05151_),
    .S(_05354_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _10213_ (.A(_05366_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(\fifo0.fifo_store[83][11] ),
    .A1(_05153_),
    .S(_05354_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _10215_ (.A(_05367_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(\fifo0.fifo_store[83][12] ),
    .A1(_05256_),
    .S(_05354_),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _10217_ (.A(_05368_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(\fifo0.fifo_store[83][13] ),
    .A1(_05211_),
    .S(_05354_),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _10219_ (.A(_05369_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(\fifo0.fifo_store[83][14] ),
    .A1(_05259_),
    .S(_05354_),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _10221_ (.A(_05370_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(\fifo0.fifo_store[83][15] ),
    .A1(_05214_),
    .S(_05354_),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _10223_ (.A(_05371_),
    .X(_01190_));
 sky130_fd_sc_hd__nor2_8 _10224_ (.A(_04052_),
    .B(_04690_),
    .Y(_05372_));
 sky130_fd_sc_hd__buf_8 _10225_ (.A(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(\fifo0.fifo_store[51][0] ),
    .A1(_05235_),
    .S(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _10227_ (.A(_05374_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _10228_ (.A0(\fifo0.fifo_store[51][1] ),
    .A1(_05198_),
    .S(_05373_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _10229_ (.A(_05375_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(\fifo0.fifo_store[51][2] ),
    .A1(_05240_),
    .S(_05373_),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _10231_ (.A(_05376_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(\fifo0.fifo_store[51][3] ),
    .A1(_05242_),
    .S(_05373_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _10233_ (.A(_05377_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\fifo0.fifo_store[51][4] ),
    .A1(_05244_),
    .S(_05373_),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_1 _10235_ (.A(_05378_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(\fifo0.fifo_store[51][5] ),
    .A1(_05144_),
    .S(_05373_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _10237_ (.A(_05379_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\fifo0.fifo_store[51][6] ),
    .A1(_05247_),
    .S(_05373_),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_1 _10239_ (.A(_05380_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(\fifo0.fifo_store[51][7] ),
    .A1(_05147_),
    .S(_05373_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _10241_ (.A(_05381_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(\fifo0.fifo_store[51][8] ),
    .A1(_05250_),
    .S(_05373_),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_1 _10243_ (.A(_05382_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(\fifo0.fifo_store[51][9] ),
    .A1(_05252_),
    .S(_05373_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _10245_ (.A(_05383_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(\fifo0.fifo_store[51][10] ),
    .A1(_05151_),
    .S(_05372_),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _10247_ (.A(_05384_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\fifo0.fifo_store[51][11] ),
    .A1(_05153_),
    .S(_05372_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _10249_ (.A(_05385_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(\fifo0.fifo_store[51][12] ),
    .A1(_05256_),
    .S(_05372_),
    .X(_05386_));
 sky130_fd_sc_hd__clkbuf_1 _10251_ (.A(_05386_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(\fifo0.fifo_store[51][13] ),
    .A1(_05211_),
    .S(_05372_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _10253_ (.A(_05387_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10254_ (.A0(\fifo0.fifo_store[51][14] ),
    .A1(_05259_),
    .S(_05372_),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _10255_ (.A(_05388_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(\fifo0.fifo_store[51][15] ),
    .A1(_05214_),
    .S(_05372_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _10257_ (.A(_05389_),
    .X(_01206_));
 sky130_fd_sc_hd__nor2_8 _10258_ (.A(_03989_),
    .B(_04297_),
    .Y(_05390_));
 sky130_fd_sc_hd__clkbuf_16 _10259_ (.A(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _10260_ (.A0(\fifo0.fifo_store[106][0] ),
    .A1(_05235_),
    .S(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _10261_ (.A(_05392_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10262_ (.A0(\fifo0.fifo_store[106][1] ),
    .A1(_05198_),
    .S(_05391_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _10263_ (.A(_05393_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(\fifo0.fifo_store[106][2] ),
    .A1(_05240_),
    .S(_05391_),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _10265_ (.A(_05394_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10266_ (.A0(\fifo0.fifo_store[106][3] ),
    .A1(_05242_),
    .S(_05391_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _10267_ (.A(_05395_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _10268_ (.A0(\fifo0.fifo_store[106][4] ),
    .A1(_05244_),
    .S(_05391_),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _10269_ (.A(_05396_),
    .X(_01211_));
 sky130_fd_sc_hd__buf_4 _10270_ (.A(_03838_),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\fifo0.fifo_store[106][5] ),
    .A1(_05397_),
    .S(_05391_),
    .X(_05398_));
 sky130_fd_sc_hd__clkbuf_1 _10272_ (.A(_05398_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\fifo0.fifo_store[106][6] ),
    .A1(_05247_),
    .S(_05391_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _10274_ (.A(_05399_),
    .X(_01213_));
 sky130_fd_sc_hd__clkbuf_4 _10275_ (.A(_03843_),
    .X(_05400_));
 sky130_fd_sc_hd__mux2_1 _10276_ (.A0(\fifo0.fifo_store[106][7] ),
    .A1(_05400_),
    .S(_05391_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _10277_ (.A(_05401_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\fifo0.fifo_store[106][8] ),
    .A1(_05250_),
    .S(_05391_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _10279_ (.A(_05402_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(\fifo0.fifo_store[106][9] ),
    .A1(_05252_),
    .S(_05391_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _10281_ (.A(_05403_),
    .X(_01216_));
 sky130_fd_sc_hd__clkbuf_4 _10282_ (.A(_03850_),
    .X(_05404_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(\fifo0.fifo_store[106][10] ),
    .A1(_05404_),
    .S(_05390_),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _10284_ (.A(_05405_),
    .X(_01217_));
 sky130_fd_sc_hd__buf_4 _10285_ (.A(_03853_),
    .X(_05406_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(\fifo0.fifo_store[106][11] ),
    .A1(_05406_),
    .S(_05390_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _10287_ (.A(_05407_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(\fifo0.fifo_store[106][12] ),
    .A1(_05256_),
    .S(_05390_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _10289_ (.A(_05408_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\fifo0.fifo_store[106][13] ),
    .A1(_05211_),
    .S(_05390_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_05409_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _10292_ (.A0(\fifo0.fifo_store[106][14] ),
    .A1(_05259_),
    .S(_05390_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _10293_ (.A(_05410_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(\fifo0.fifo_store[106][15] ),
    .A1(_05214_),
    .S(_05390_),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _10295_ (.A(_05411_),
    .X(_01222_));
 sky130_fd_sc_hd__nor2_8 _10296_ (.A(_03868_),
    .B(_03990_),
    .Y(_05412_));
 sky130_fd_sc_hd__buf_6 _10297_ (.A(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(\fifo0.fifo_store[82][0] ),
    .A1(_05235_),
    .S(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_1 _10299_ (.A(_05414_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10300_ (.A0(\fifo0.fifo_store[82][1] ),
    .A1(_05198_),
    .S(_05413_),
    .X(_05415_));
 sky130_fd_sc_hd__clkbuf_1 _10301_ (.A(_05415_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(\fifo0.fifo_store[82][2] ),
    .A1(_05240_),
    .S(_05413_),
    .X(_05416_));
 sky130_fd_sc_hd__clkbuf_1 _10303_ (.A(_05416_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(\fifo0.fifo_store[82][3] ),
    .A1(_05242_),
    .S(_05413_),
    .X(_05417_));
 sky130_fd_sc_hd__clkbuf_1 _10305_ (.A(_05417_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10306_ (.A0(\fifo0.fifo_store[82][4] ),
    .A1(_05244_),
    .S(_05413_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _10307_ (.A(_05418_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10308_ (.A0(\fifo0.fifo_store[82][5] ),
    .A1(_05397_),
    .S(_05413_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _10309_ (.A(_05419_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _10310_ (.A0(\fifo0.fifo_store[82][6] ),
    .A1(_05247_),
    .S(_05413_),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _10311_ (.A(_05420_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(\fifo0.fifo_store[82][7] ),
    .A1(_05400_),
    .S(_05413_),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _10313_ (.A(_05421_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\fifo0.fifo_store[82][8] ),
    .A1(_05250_),
    .S(_05413_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _10315_ (.A(_05422_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\fifo0.fifo_store[82][9] ),
    .A1(_05252_),
    .S(_05413_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _10317_ (.A(_05423_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\fifo0.fifo_store[82][10] ),
    .A1(_05404_),
    .S(_05412_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_05424_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\fifo0.fifo_store[82][11] ),
    .A1(_05406_),
    .S(_05412_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _10321_ (.A(_05425_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\fifo0.fifo_store[82][12] ),
    .A1(_05256_),
    .S(_05412_),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_1 _10323_ (.A(_05426_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\fifo0.fifo_store[82][13] ),
    .A1(_05211_),
    .S(_05412_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_1 _10325_ (.A(_05427_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(\fifo0.fifo_store[82][14] ),
    .A1(_05259_),
    .S(_05412_),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_1 _10327_ (.A(_05428_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(\fifo0.fifo_store[82][15] ),
    .A1(_05214_),
    .S(_05412_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _10329_ (.A(_05429_),
    .X(_01238_));
 sky130_fd_sc_hd__nor2_8 _10330_ (.A(_03868_),
    .B(_04032_),
    .Y(_05430_));
 sky130_fd_sc_hd__buf_6 _10331_ (.A(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(\fifo0.fifo_store[81][0] ),
    .A1(_05235_),
    .S(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _10333_ (.A(_05432_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(\fifo0.fifo_store[81][1] ),
    .A1(_05198_),
    .S(_05431_),
    .X(_05433_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(_05433_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\fifo0.fifo_store[81][2] ),
    .A1(_05240_),
    .S(_05431_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_1 _10337_ (.A(_05434_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(\fifo0.fifo_store[81][3] ),
    .A1(_05242_),
    .S(_05431_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _10339_ (.A(_05435_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _10340_ (.A0(\fifo0.fifo_store[81][4] ),
    .A1(_05244_),
    .S(_05431_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _10341_ (.A(_05436_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\fifo0.fifo_store[81][5] ),
    .A1(_05397_),
    .S(_05431_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _10343_ (.A(_05437_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\fifo0.fifo_store[81][6] ),
    .A1(_05247_),
    .S(_05431_),
    .X(_05438_));
 sky130_fd_sc_hd__clkbuf_1 _10345_ (.A(_05438_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(\fifo0.fifo_store[81][7] ),
    .A1(_05400_),
    .S(_05431_),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_1 _10347_ (.A(_05439_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(\fifo0.fifo_store[81][8] ),
    .A1(_05250_),
    .S(_05431_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _10349_ (.A(_05440_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _10350_ (.A0(\fifo0.fifo_store[81][9] ),
    .A1(_05252_),
    .S(_05431_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_1 _10351_ (.A(_05441_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _10352_ (.A0(\fifo0.fifo_store[81][10] ),
    .A1(_05404_),
    .S(_05430_),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _10353_ (.A(_05442_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(\fifo0.fifo_store[81][11] ),
    .A1(_05406_),
    .S(_05430_),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_1 _10355_ (.A(_05443_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _10356_ (.A0(\fifo0.fifo_store[81][12] ),
    .A1(_05256_),
    .S(_05430_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _10357_ (.A(_05444_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10358_ (.A0(\fifo0.fifo_store[81][13] ),
    .A1(_05211_),
    .S(_05430_),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_1 _10359_ (.A(_05445_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10360_ (.A0(\fifo0.fifo_store[81][14] ),
    .A1(_05259_),
    .S(_05430_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _10361_ (.A(_05446_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(\fifo0.fifo_store[81][15] ),
    .A1(_05214_),
    .S(_05430_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_1 _10363_ (.A(_05447_),
    .X(_01254_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(_04201_),
    .B(_04172_),
    .X(_05448_));
 sky130_fd_sc_hd__buf_4 _10365_ (.A(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__clkbuf_16 _10366_ (.A(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[94][0] ),
    .S(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _10368_ (.A(_05451_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[94][1] ),
    .S(_05450_),
    .X(_05452_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_05452_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[94][2] ),
    .S(_05450_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _10372_ (.A(_05453_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[94][3] ),
    .S(_05450_),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_05454_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[94][4] ),
    .S(_05450_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_1 _10376_ (.A(_05455_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _10377_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[94][5] ),
    .S(_05450_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _10378_ (.A(_05456_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _10379_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[94][6] ),
    .S(_05450_),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _10380_ (.A(_05457_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _10381_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[94][7] ),
    .S(_05450_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(_05458_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[94][8] ),
    .S(_05450_),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_1 _10384_ (.A(_05459_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[94][9] ),
    .S(_05450_),
    .X(_05460_));
 sky130_fd_sc_hd__clkbuf_1 _10386_ (.A(_05460_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _10387_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[94][10] ),
    .S(_05449_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _10388_ (.A(_05461_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _10389_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[94][11] ),
    .S(_05449_),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_1 _10390_ (.A(_05462_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _10391_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[94][12] ),
    .S(_05449_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _10392_ (.A(_05463_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _10393_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[94][13] ),
    .S(_05449_),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_1 _10394_ (.A(_05464_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[94][14] ),
    .S(_05449_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _10396_ (.A(_05465_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[94][15] ),
    .S(_05449_),
    .X(_05466_));
 sky130_fd_sc_hd__clkbuf_1 _10398_ (.A(_05466_),
    .X(_01270_));
 sky130_fd_sc_hd__nor2_8 _10399_ (.A(_04277_),
    .B(_04629_),
    .Y(_05467_));
 sky130_fd_sc_hd__buf_6 _10400_ (.A(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(\fifo0.fifo_store[44][0] ),
    .A1(_05235_),
    .S(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__clkbuf_1 _10402_ (.A(_05469_),
    .X(_01271_));
 sky130_fd_sc_hd__buf_4 _10403_ (.A(_03872_),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(\fifo0.fifo_store[44][1] ),
    .A1(_05470_),
    .S(_05468_),
    .X(_05471_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_05471_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(\fifo0.fifo_store[44][2] ),
    .A1(_05240_),
    .S(_05468_),
    .X(_05472_));
 sky130_fd_sc_hd__clkbuf_1 _10407_ (.A(_05472_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(\fifo0.fifo_store[44][3] ),
    .A1(_05242_),
    .S(_05468_),
    .X(_05473_));
 sky130_fd_sc_hd__clkbuf_1 _10409_ (.A(_05473_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(\fifo0.fifo_store[44][4] ),
    .A1(_05244_),
    .S(_05468_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _10411_ (.A(_05474_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(\fifo0.fifo_store[44][5] ),
    .A1(_05397_),
    .S(_05468_),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _10413_ (.A(_05475_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(\fifo0.fifo_store[44][6] ),
    .A1(_05247_),
    .S(_05468_),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_05476_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(\fifo0.fifo_store[44][7] ),
    .A1(_05400_),
    .S(_05468_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_05477_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\fifo0.fifo_store[44][8] ),
    .A1(_05250_),
    .S(_05468_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_05478_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\fifo0.fifo_store[44][9] ),
    .A1(_05252_),
    .S(_05468_),
    .X(_05479_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_05479_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\fifo0.fifo_store[44][10] ),
    .A1(_05404_),
    .S(_05467_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_05480_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\fifo0.fifo_store[44][11] ),
    .A1(_05406_),
    .S(_05467_),
    .X(_05481_));
 sky130_fd_sc_hd__clkbuf_1 _10425_ (.A(_05481_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\fifo0.fifo_store[44][12] ),
    .A1(_05256_),
    .S(_05467_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_05482_),
    .X(_01283_));
 sky130_fd_sc_hd__clkbuf_4 _10428_ (.A(_03908_),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _10429_ (.A0(\fifo0.fifo_store[44][13] ),
    .A1(_05483_),
    .S(_05467_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_05484_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(\fifo0.fifo_store[44][14] ),
    .A1(_05259_),
    .S(_05467_),
    .X(_05485_));
 sky130_fd_sc_hd__clkbuf_1 _10432_ (.A(_05485_),
    .X(_01285_));
 sky130_fd_sc_hd__buf_2 _10433_ (.A(_03914_),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_1 _10434_ (.A0(\fifo0.fifo_store[44][15] ),
    .A1(_05486_),
    .S(_05467_),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_1 _10435_ (.A(_05487_),
    .X(_01286_));
 sky130_fd_sc_hd__buf_4 _10436_ (.A(_03821_),
    .X(_05488_));
 sky130_fd_sc_hd__nor2_8 _10437_ (.A(_04052_),
    .B(_04629_),
    .Y(_05489_));
 sky130_fd_sc_hd__buf_8 _10438_ (.A(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(\fifo0.fifo_store[43][0] ),
    .A1(_05488_),
    .S(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_05491_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\fifo0.fifo_store[43][1] ),
    .A1(_05470_),
    .S(_05490_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_05492_),
    .X(_01288_));
 sky130_fd_sc_hd__clkbuf_4 _10443_ (.A(_03875_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _10444_ (.A0(\fifo0.fifo_store[43][2] ),
    .A1(_05493_),
    .S(_05490_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _10445_ (.A(_05494_),
    .X(_01289_));
 sky130_fd_sc_hd__buf_2 _10446_ (.A(_03878_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(\fifo0.fifo_store[43][3] ),
    .A1(_05495_),
    .S(_05490_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _10448_ (.A(_05496_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _10449_ (.A(_03881_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(\fifo0.fifo_store[43][4] ),
    .A1(_05497_),
    .S(_05490_),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _10451_ (.A(_05498_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(\fifo0.fifo_store[43][5] ),
    .A1(_05397_),
    .S(_05490_),
    .X(_05499_));
 sky130_fd_sc_hd__clkbuf_1 _10453_ (.A(_05499_),
    .X(_01292_));
 sky130_fd_sc_hd__clkbuf_4 _10454_ (.A(_03887_),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(\fifo0.fifo_store[43][6] ),
    .A1(_05500_),
    .S(_05490_),
    .X(_05501_));
 sky130_fd_sc_hd__clkbuf_1 _10456_ (.A(_05501_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(\fifo0.fifo_store[43][7] ),
    .A1(_05400_),
    .S(_05490_),
    .X(_05502_));
 sky130_fd_sc_hd__clkbuf_1 _10458_ (.A(_05502_),
    .X(_01294_));
 sky130_fd_sc_hd__clkbuf_4 _10459_ (.A(_03893_),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\fifo0.fifo_store[43][8] ),
    .A1(_05503_),
    .S(_05490_),
    .X(_05504_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_05504_),
    .X(_01295_));
 sky130_fd_sc_hd__buf_2 _10462_ (.A(_03896_),
    .X(_05505_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(\fifo0.fifo_store[43][9] ),
    .A1(_05505_),
    .S(_05490_),
    .X(_05506_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(_05506_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(\fifo0.fifo_store[43][10] ),
    .A1(_05404_),
    .S(_05489_),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _10466_ (.A(_05507_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(\fifo0.fifo_store[43][11] ),
    .A1(_05406_),
    .S(_05489_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(_05508_),
    .X(_01298_));
 sky130_fd_sc_hd__buf_4 _10469_ (.A(_03905_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(\fifo0.fifo_store[43][12] ),
    .A1(_05509_),
    .S(_05489_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_1 _10471_ (.A(_05510_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\fifo0.fifo_store[43][13] ),
    .A1(_05483_),
    .S(_05489_),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(_05511_),
    .X(_01300_));
 sky130_fd_sc_hd__buf_4 _10474_ (.A(_03911_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(\fifo0.fifo_store[43][14] ),
    .A1(_05512_),
    .S(_05489_),
    .X(_05513_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_05513_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\fifo0.fifo_store[43][15] ),
    .A1(_05486_),
    .S(_05489_),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_05514_),
    .X(_01302_));
 sky130_fd_sc_hd__nor2_8 _10479_ (.A(_03989_),
    .B(_04629_),
    .Y(_05515_));
 sky130_fd_sc_hd__buf_8 _10480_ (.A(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(\fifo0.fifo_store[42][0] ),
    .A1(_05488_),
    .S(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_05517_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\fifo0.fifo_store[42][1] ),
    .A1(_05470_),
    .S(_05516_),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_05518_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\fifo0.fifo_store[42][2] ),
    .A1(_05493_),
    .S(_05516_),
    .X(_05519_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_05519_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\fifo0.fifo_store[42][3] ),
    .A1(_05495_),
    .S(_05516_),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_05520_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\fifo0.fifo_store[42][4] ),
    .A1(_05497_),
    .S(_05516_),
    .X(_05521_));
 sky130_fd_sc_hd__clkbuf_1 _10490_ (.A(_05521_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\fifo0.fifo_store[42][5] ),
    .A1(_05397_),
    .S(_05516_),
    .X(_05522_));
 sky130_fd_sc_hd__clkbuf_1 _10492_ (.A(_05522_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(\fifo0.fifo_store[42][6] ),
    .A1(_05500_),
    .S(_05516_),
    .X(_05523_));
 sky130_fd_sc_hd__clkbuf_1 _10494_ (.A(_05523_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\fifo0.fifo_store[42][7] ),
    .A1(_05400_),
    .S(_05516_),
    .X(_05524_));
 sky130_fd_sc_hd__clkbuf_1 _10496_ (.A(_05524_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(\fifo0.fifo_store[42][8] ),
    .A1(_05503_),
    .S(_05516_),
    .X(_05525_));
 sky130_fd_sc_hd__clkbuf_1 _10498_ (.A(_05525_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(\fifo0.fifo_store[42][9] ),
    .A1(_05505_),
    .S(_05516_),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_1 _10500_ (.A(_05526_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\fifo0.fifo_store[42][10] ),
    .A1(_05404_),
    .S(_05515_),
    .X(_05527_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_05527_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(\fifo0.fifo_store[42][11] ),
    .A1(_05406_),
    .S(_05515_),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _10504_ (.A(_05528_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(\fifo0.fifo_store[42][12] ),
    .A1(_05509_),
    .S(_05515_),
    .X(_05529_));
 sky130_fd_sc_hd__clkbuf_1 _10506_ (.A(_05529_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\fifo0.fifo_store[42][13] ),
    .A1(_05483_),
    .S(_05515_),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(_05530_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(\fifo0.fifo_store[42][14] ),
    .A1(_05512_),
    .S(_05515_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_05531_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\fifo0.fifo_store[42][15] ),
    .A1(_05486_),
    .S(_05515_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(_05532_),
    .X(_01318_));
 sky130_fd_sc_hd__nor2_4 _10513_ (.A(_04031_),
    .B(_04629_),
    .Y(_05533_));
 sky130_fd_sc_hd__buf_8 _10514_ (.A(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\fifo0.fifo_store[41][0] ),
    .A1(_05488_),
    .S(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_05535_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\fifo0.fifo_store[41][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_05534_),
    .X(_05536_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_05536_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\fifo0.fifo_store[41][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_05534_),
    .X(_05537_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_05537_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\fifo0.fifo_store[41][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_05534_),
    .X(_05538_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_05538_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(\fifo0.fifo_store[41][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_05534_),
    .X(_05539_));
 sky130_fd_sc_hd__clkbuf_1 _10524_ (.A(_05539_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\fifo0.fifo_store[41][5] ),
    .A1(_05397_),
    .S(_05534_),
    .X(_05540_));
 sky130_fd_sc_hd__clkbuf_1 _10526_ (.A(_05540_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\fifo0.fifo_store[41][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_05534_),
    .X(_05541_));
 sky130_fd_sc_hd__clkbuf_1 _10528_ (.A(_05541_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\fifo0.fifo_store[41][7] ),
    .A1(_05400_),
    .S(_05534_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _10530_ (.A(_05542_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\fifo0.fifo_store[41][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_05534_),
    .X(_05543_));
 sky130_fd_sc_hd__clkbuf_1 _10532_ (.A(_05543_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\fifo0.fifo_store[41][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_05534_),
    .X(_05544_));
 sky130_fd_sc_hd__clkbuf_1 _10534_ (.A(_05544_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(\fifo0.fifo_store[41][10] ),
    .A1(_05404_),
    .S(_05533_),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _10536_ (.A(_05545_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(\fifo0.fifo_store[41][11] ),
    .A1(_05406_),
    .S(_05533_),
    .X(_05546_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(_05546_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\fifo0.fifo_store[41][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_05533_),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(_05547_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\fifo0.fifo_store[41][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_05533_),
    .X(_05548_));
 sky130_fd_sc_hd__clkbuf_1 _10542_ (.A(_05548_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(\fifo0.fifo_store[41][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_05533_),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(_05549_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(\fifo0.fifo_store[41][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_05533_),
    .X(_05550_));
 sky130_fd_sc_hd__clkbuf_1 _10546_ (.A(_05550_),
    .X(_01334_));
 sky130_fd_sc_hd__nor2_4 _10547_ (.A(_03815_),
    .B(_04629_),
    .Y(_05551_));
 sky130_fd_sc_hd__buf_8 _10548_ (.A(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_1 _10549_ (.A0(\fifo0.fifo_store[40][0] ),
    .A1(_05488_),
    .S(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__clkbuf_1 _10550_ (.A(_05553_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(\fifo0.fifo_store[40][1] ),
    .A1(_05470_),
    .S(_05552_),
    .X(_05554_));
 sky130_fd_sc_hd__clkbuf_1 _10552_ (.A(_05554_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(\fifo0.fifo_store[40][2] ),
    .A1(_05493_),
    .S(_05552_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _10554_ (.A(_05555_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\fifo0.fifo_store[40][3] ),
    .A1(_05495_),
    .S(_05552_),
    .X(_05556_));
 sky130_fd_sc_hd__clkbuf_1 _10556_ (.A(_05556_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(\fifo0.fifo_store[40][4] ),
    .A1(_05497_),
    .S(_05552_),
    .X(_05557_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_05557_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\fifo0.fifo_store[40][5] ),
    .A1(_05397_),
    .S(_05552_),
    .X(_05558_));
 sky130_fd_sc_hd__clkbuf_1 _10560_ (.A(_05558_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(\fifo0.fifo_store[40][6] ),
    .A1(_05500_),
    .S(_05552_),
    .X(_05559_));
 sky130_fd_sc_hd__clkbuf_1 _10562_ (.A(_05559_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(\fifo0.fifo_store[40][7] ),
    .A1(_05400_),
    .S(_05552_),
    .X(_05560_));
 sky130_fd_sc_hd__clkbuf_1 _10564_ (.A(_05560_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10565_ (.A0(\fifo0.fifo_store[40][8] ),
    .A1(_05503_),
    .S(_05552_),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _10566_ (.A(_05561_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\fifo0.fifo_store[40][9] ),
    .A1(_05505_),
    .S(_05552_),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_05562_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(\fifo0.fifo_store[40][10] ),
    .A1(_05404_),
    .S(_05551_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_05563_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(\fifo0.fifo_store[40][11] ),
    .A1(_05406_),
    .S(_05551_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_05564_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\fifo0.fifo_store[40][12] ),
    .A1(_05509_),
    .S(_05551_),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_05565_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\fifo0.fifo_store[40][13] ),
    .A1(_05483_),
    .S(_05551_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _10576_ (.A(_05566_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(\fifo0.fifo_store[40][14] ),
    .A1(_05512_),
    .S(_05551_),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _10578_ (.A(_05567_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(\fifo0.fifo_store[40][15] ),
    .A1(_05486_),
    .S(_05551_),
    .X(_05568_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(_05568_),
    .X(_01350_));
 sky130_fd_sc_hd__nor2_8 _10581_ (.A(_03814_),
    .B(_04053_),
    .Y(_05569_));
 sky130_fd_sc_hd__buf_6 _10582_ (.A(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\fifo0.fifo_store[3][0] ),
    .A1(_05488_),
    .S(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_05571_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\fifo0.fifo_store[3][1] ),
    .A1(_05470_),
    .S(_05570_),
    .X(_05572_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_05572_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(\fifo0.fifo_store[3][2] ),
    .A1(_05493_),
    .S(_05570_),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _10588_ (.A(_05573_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\fifo0.fifo_store[3][3] ),
    .A1(_05495_),
    .S(_05570_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(_05574_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\fifo0.fifo_store[3][4] ),
    .A1(_05497_),
    .S(_05570_),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _10592_ (.A(_05575_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(\fifo0.fifo_store[3][5] ),
    .A1(_05397_),
    .S(_05570_),
    .X(_05576_));
 sky130_fd_sc_hd__clkbuf_1 _10594_ (.A(_05576_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(\fifo0.fifo_store[3][6] ),
    .A1(_05500_),
    .S(_05570_),
    .X(_05577_));
 sky130_fd_sc_hd__clkbuf_1 _10596_ (.A(_05577_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\fifo0.fifo_store[3][7] ),
    .A1(_05400_),
    .S(_05570_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _10598_ (.A(_05578_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(\fifo0.fifo_store[3][8] ),
    .A1(_05503_),
    .S(_05570_),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(_05579_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\fifo0.fifo_store[3][9] ),
    .A1(_05505_),
    .S(_05570_),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_05580_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\fifo0.fifo_store[3][10] ),
    .A1(_05404_),
    .S(_05569_),
    .X(_05581_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_05581_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\fifo0.fifo_store[3][11] ),
    .A1(_05406_),
    .S(_05569_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_05582_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\fifo0.fifo_store[3][12] ),
    .A1(_05509_),
    .S(_05569_),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_05583_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\fifo0.fifo_store[3][13] ),
    .A1(_05483_),
    .S(_05569_),
    .X(_05584_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_05584_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\fifo0.fifo_store[3][14] ),
    .A1(_05512_),
    .S(_05569_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_05585_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\fifo0.fifo_store[3][15] ),
    .A1(_05486_),
    .S(_05569_),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_05586_),
    .X(_01366_));
 sky130_fd_sc_hd__or2_1 _10615_ (.A(_03806_),
    .B(_04627_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_8 _10616_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__or2_1 _10617_ (.A(_04201_),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_4 _10618_ (.A(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__buf_8 _10619_ (.A(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[38][0] ),
    .S(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_05592_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[38][1] ),
    .S(_05591_),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_05593_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[38][2] ),
    .S(_05591_),
    .X(_05594_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_05594_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[38][3] ),
    .S(_05591_),
    .X(_05595_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_05595_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[38][4] ),
    .S(_05591_),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_05596_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[38][5] ),
    .S(_05591_),
    .X(_05597_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_05597_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[38][6] ),
    .S(_05591_),
    .X(_05598_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_05598_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[38][7] ),
    .S(_05591_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_05599_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[38][8] ),
    .S(_05591_),
    .X(_05600_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_05600_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[38][9] ),
    .S(_05591_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_05601_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[38][10] ),
    .S(_05590_),
    .X(_05602_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_05602_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[38][11] ),
    .S(_05590_),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_1 _10643_ (.A(_05603_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[38][12] ),
    .S(_05590_),
    .X(_05604_));
 sky130_fd_sc_hd__clkbuf_1 _10645_ (.A(_05604_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[38][13] ),
    .S(_05590_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_1 _10647_ (.A(_05605_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[38][14] ),
    .S(_05590_),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_1 _10649_ (.A(_05606_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[38][15] ),
    .S(_05590_),
    .X(_05607_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_05607_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_8 _10652_ (.A(_03964_),
    .B(_05588_),
    .Y(_05608_));
 sky130_fd_sc_hd__buf_6 _10653_ (.A(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(\fifo0.fifo_store[37][0] ),
    .A1(_05488_),
    .S(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(_05610_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\fifo0.fifo_store[37][1] ),
    .A1(_05470_),
    .S(_05609_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(_05611_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(\fifo0.fifo_store[37][2] ),
    .A1(_05493_),
    .S(_05609_),
    .X(_05612_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(_05612_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\fifo0.fifo_store[37][3] ),
    .A1(_05495_),
    .S(_05609_),
    .X(_05613_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(_05613_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\fifo0.fifo_store[37][4] ),
    .A1(_05497_),
    .S(_05609_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_05614_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\fifo0.fifo_store[37][5] ),
    .A1(_05397_),
    .S(_05609_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_05615_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\fifo0.fifo_store[37][6] ),
    .A1(_05500_),
    .S(_05609_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_05616_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\fifo0.fifo_store[37][7] ),
    .A1(_05400_),
    .S(_05609_),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_05617_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\fifo0.fifo_store[37][8] ),
    .A1(_05503_),
    .S(_05609_),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_05618_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\fifo0.fifo_store[37][9] ),
    .A1(_05505_),
    .S(_05609_),
    .X(_05619_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_05619_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\fifo0.fifo_store[37][10] ),
    .A1(_05404_),
    .S(_05608_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_05620_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\fifo0.fifo_store[37][11] ),
    .A1(_05406_),
    .S(_05608_),
    .X(_05621_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_05621_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\fifo0.fifo_store[37][12] ),
    .A1(_05509_),
    .S(_05608_),
    .X(_05622_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_05622_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\fifo0.fifo_store[37][13] ),
    .A1(_05483_),
    .S(_05608_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_05623_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\fifo0.fifo_store[37][14] ),
    .A1(_05512_),
    .S(_05608_),
    .X(_05624_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_05624_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\fifo0.fifo_store[37][15] ),
    .A1(_05486_),
    .S(_05608_),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_1 _10685_ (.A(_05625_),
    .X(_01398_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(_03943_),
    .B(_04356_),
    .X(_05626_));
 sky130_fd_sc_hd__buf_4 _10687_ (.A(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__buf_8 _10688_ (.A(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[14][0] ),
    .S(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(_05629_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[14][1] ),
    .S(_05628_),
    .X(_05630_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(_05630_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[14][2] ),
    .S(_05628_),
    .X(_05631_));
 sky130_fd_sc_hd__clkbuf_1 _10694_ (.A(_05631_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[14][3] ),
    .S(_05628_),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_05632_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[14][4] ),
    .S(_05628_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_1 _10698_ (.A(_05633_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[14][5] ),
    .S(_05628_),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_05634_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[14][6] ),
    .S(_05628_),
    .X(_05635_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_05635_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[14][7] ),
    .S(_05628_),
    .X(_05636_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_05636_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[14][8] ),
    .S(_05628_),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _10706_ (.A(_05637_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[14][9] ),
    .S(_05628_),
    .X(_05638_));
 sky130_fd_sc_hd__clkbuf_1 _10708_ (.A(_05638_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[14][10] ),
    .S(_05627_),
    .X(_05639_));
 sky130_fd_sc_hd__clkbuf_1 _10710_ (.A(_05639_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[14][11] ),
    .S(_05627_),
    .X(_05640_));
 sky130_fd_sc_hd__clkbuf_1 _10712_ (.A(_05640_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[14][12] ),
    .S(_05627_),
    .X(_05641_));
 sky130_fd_sc_hd__clkbuf_1 _10714_ (.A(_05641_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[14][13] ),
    .S(_05627_),
    .X(_05642_));
 sky130_fd_sc_hd__clkbuf_1 _10716_ (.A(_05642_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[14][14] ),
    .S(_05627_),
    .X(_05643_));
 sky130_fd_sc_hd__clkbuf_1 _10718_ (.A(_05643_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[14][15] ),
    .S(_05627_),
    .X(_05644_));
 sky130_fd_sc_hd__clkbuf_1 _10720_ (.A(_05644_),
    .X(_01414_));
 sky130_fd_sc_hd__nor2_8 _10721_ (.A(_04277_),
    .B(_05588_),
    .Y(_05645_));
 sky130_fd_sc_hd__buf_6 _10722_ (.A(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(\fifo0.fifo_store[36][0] ),
    .A1(_05488_),
    .S(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(_05647_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\fifo0.fifo_store[36][1] ),
    .A1(_05470_),
    .S(_05646_),
    .X(_05648_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_05648_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(\fifo0.fifo_store[36][2] ),
    .A1(_05493_),
    .S(_05646_),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_05649_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(\fifo0.fifo_store[36][3] ),
    .A1(_05495_),
    .S(_05646_),
    .X(_05650_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_05650_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(\fifo0.fifo_store[36][4] ),
    .A1(_05497_),
    .S(_05646_),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(_05651_),
    .X(_01419_));
 sky130_fd_sc_hd__clkbuf_8 _10733_ (.A(_03838_),
    .X(_05652_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\fifo0.fifo_store[36][5] ),
    .A1(_05652_),
    .S(_05646_),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_05653_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\fifo0.fifo_store[36][6] ),
    .A1(_05500_),
    .S(_05646_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_05654_),
    .X(_01421_));
 sky130_fd_sc_hd__buf_4 _10738_ (.A(_03843_),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\fifo0.fifo_store[36][7] ),
    .A1(_05655_),
    .S(_05646_),
    .X(_05656_));
 sky130_fd_sc_hd__clkbuf_1 _10740_ (.A(_05656_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\fifo0.fifo_store[36][8] ),
    .A1(_05503_),
    .S(_05646_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_1 _10742_ (.A(_05657_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\fifo0.fifo_store[36][9] ),
    .A1(_05505_),
    .S(_05646_),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_05658_),
    .X(_01424_));
 sky130_fd_sc_hd__buf_4 _10745_ (.A(_03850_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\fifo0.fifo_store[36][10] ),
    .A1(_05659_),
    .S(_05645_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_05660_),
    .X(_01425_));
 sky130_fd_sc_hd__buf_6 _10748_ (.A(_03853_),
    .X(_05661_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\fifo0.fifo_store[36][11] ),
    .A1(_05661_),
    .S(_05645_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _10750_ (.A(_05662_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\fifo0.fifo_store[36][12] ),
    .A1(_05509_),
    .S(_05645_),
    .X(_05663_));
 sky130_fd_sc_hd__clkbuf_1 _10752_ (.A(_05663_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\fifo0.fifo_store[36][13] ),
    .A1(_05483_),
    .S(_05645_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_1 _10754_ (.A(_05664_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(\fifo0.fifo_store[36][14] ),
    .A1(_05512_),
    .S(_05645_),
    .X(_05665_));
 sky130_fd_sc_hd__clkbuf_1 _10756_ (.A(_05665_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(\fifo0.fifo_store[36][15] ),
    .A1(_05486_),
    .S(_05645_),
    .X(_05666_));
 sky130_fd_sc_hd__clkbuf_1 _10758_ (.A(_05666_),
    .X(_01430_));
 sky130_fd_sc_hd__nor2_4 _10759_ (.A(_04052_),
    .B(_05588_),
    .Y(_05667_));
 sky130_fd_sc_hd__buf_6 _10760_ (.A(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(\fifo0.fifo_store[35][0] ),
    .A1(_05488_),
    .S(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__clkbuf_1 _10762_ (.A(_05669_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(\fifo0.fifo_store[35][1] ),
    .A1(_05470_),
    .S(_05668_),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_1 _10764_ (.A(_05670_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(\fifo0.fifo_store[35][2] ),
    .A1(_05493_),
    .S(_05668_),
    .X(_05671_));
 sky130_fd_sc_hd__clkbuf_1 _10766_ (.A(_05671_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(\fifo0.fifo_store[35][3] ),
    .A1(_05495_),
    .S(_05668_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _10768_ (.A(_05672_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(\fifo0.fifo_store[35][4] ),
    .A1(_05497_),
    .S(_05668_),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_1 _10770_ (.A(_05673_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\fifo0.fifo_store[35][5] ),
    .A1(_05652_),
    .S(_05668_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _10772_ (.A(_05674_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\fifo0.fifo_store[35][6] ),
    .A1(_05500_),
    .S(_05668_),
    .X(_05675_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_05675_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\fifo0.fifo_store[35][7] ),
    .A1(_05655_),
    .S(_05668_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_05676_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\fifo0.fifo_store[35][8] ),
    .A1(_05503_),
    .S(_05668_),
    .X(_05677_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_05677_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\fifo0.fifo_store[35][9] ),
    .A1(_05505_),
    .S(_05668_),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_05678_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\fifo0.fifo_store[35][10] ),
    .A1(_05659_),
    .S(_05667_),
    .X(_05679_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_05679_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\fifo0.fifo_store[35][11] ),
    .A1(_05661_),
    .S(_05667_),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_05680_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\fifo0.fifo_store[35][12] ),
    .A1(_05509_),
    .S(_05667_),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_05681_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\fifo0.fifo_store[35][13] ),
    .A1(_05483_),
    .S(_05667_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_05682_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\fifo0.fifo_store[35][14] ),
    .A1(_05512_),
    .S(_05667_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_05683_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\fifo0.fifo_store[35][15] ),
    .A1(_05486_),
    .S(_05667_),
    .X(_05684_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_05684_),
    .X(_01446_));
 sky130_fd_sc_hd__nor2_4 _10793_ (.A(_03989_),
    .B(_05588_),
    .Y(_05685_));
 sky130_fd_sc_hd__buf_6 _10794_ (.A(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\fifo0.fifo_store[34][0] ),
    .A1(_05488_),
    .S(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_05687_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\fifo0.fifo_store[34][1] ),
    .A1(_05470_),
    .S(_05686_),
    .X(_05688_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_05688_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\fifo0.fifo_store[34][2] ),
    .A1(_05493_),
    .S(_05686_),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _10800_ (.A(_05689_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(\fifo0.fifo_store[34][3] ),
    .A1(_05495_),
    .S(_05686_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_05690_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(\fifo0.fifo_store[34][4] ),
    .A1(_05497_),
    .S(_05686_),
    .X(_05691_));
 sky130_fd_sc_hd__clkbuf_1 _10804_ (.A(_05691_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(\fifo0.fifo_store[34][5] ),
    .A1(_05652_),
    .S(_05686_),
    .X(_05692_));
 sky130_fd_sc_hd__clkbuf_1 _10806_ (.A(_05692_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\fifo0.fifo_store[34][6] ),
    .A1(_05500_),
    .S(_05686_),
    .X(_05693_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_05693_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(\fifo0.fifo_store[34][7] ),
    .A1(_05655_),
    .S(_05686_),
    .X(_05694_));
 sky130_fd_sc_hd__clkbuf_1 _10810_ (.A(_05694_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\fifo0.fifo_store[34][8] ),
    .A1(_05503_),
    .S(_05686_),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_1 _10812_ (.A(_05695_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(\fifo0.fifo_store[34][9] ),
    .A1(_05505_),
    .S(_05686_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_1 _10814_ (.A(_05696_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\fifo0.fifo_store[34][10] ),
    .A1(_05659_),
    .S(_05685_),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(_05697_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(\fifo0.fifo_store[34][11] ),
    .A1(_05661_),
    .S(_05685_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _10818_ (.A(_05698_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(\fifo0.fifo_store[34][12] ),
    .A1(_05509_),
    .S(_05685_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(_05699_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\fifo0.fifo_store[34][13] ),
    .A1(_05483_),
    .S(_05685_),
    .X(_05700_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_05700_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\fifo0.fifo_store[34][14] ),
    .A1(_05512_),
    .S(_05685_),
    .X(_05701_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_05701_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\fifo0.fifo_store[34][15] ),
    .A1(_05486_),
    .S(_05685_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_05702_),
    .X(_01462_));
 sky130_fd_sc_hd__nor2_8 _10827_ (.A(_03986_),
    .B(_04053_),
    .Y(_05703_));
 sky130_fd_sc_hd__buf_6 _10828_ (.A(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\fifo0.fifo_store[99][0] ),
    .A1(_05488_),
    .S(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_05705_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\fifo0.fifo_store[99][1] ),
    .A1(_05470_),
    .S(_05704_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_05706_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\fifo0.fifo_store[99][2] ),
    .A1(_05493_),
    .S(_05704_),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_05707_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\fifo0.fifo_store[99][3] ),
    .A1(_05495_),
    .S(_05704_),
    .X(_05708_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_05708_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\fifo0.fifo_store[99][4] ),
    .A1(_05497_),
    .S(_05704_),
    .X(_05709_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_05709_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\fifo0.fifo_store[99][5] ),
    .A1(_05652_),
    .S(_05704_),
    .X(_05710_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_05710_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\fifo0.fifo_store[99][6] ),
    .A1(_05500_),
    .S(_05704_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _10842_ (.A(_05711_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\fifo0.fifo_store[99][7] ),
    .A1(_05655_),
    .S(_05704_),
    .X(_05712_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_05712_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\fifo0.fifo_store[99][8] ),
    .A1(_05503_),
    .S(_05704_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_05713_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\fifo0.fifo_store[99][9] ),
    .A1(_05505_),
    .S(_05704_),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_05714_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\fifo0.fifo_store[99][10] ),
    .A1(_05659_),
    .S(_05703_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_05715_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\fifo0.fifo_store[99][11] ),
    .A1(_05661_),
    .S(_05703_),
    .X(_05716_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_05716_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\fifo0.fifo_store[99][12] ),
    .A1(_05509_),
    .S(_05703_),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_05717_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\fifo0.fifo_store[99][13] ),
    .A1(_05483_),
    .S(_05703_),
    .X(_05718_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_05718_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\fifo0.fifo_store[99][14] ),
    .A1(_05512_),
    .S(_05703_),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_05719_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\fifo0.fifo_store[99][15] ),
    .A1(_05486_),
    .S(_05703_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_05720_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_4 _10861_ (.A(_03821_),
    .X(_05721_));
 sky130_fd_sc_hd__nor2_4 _10862_ (.A(_04031_),
    .B(_05588_),
    .Y(_05722_));
 sky130_fd_sc_hd__buf_6 _10863_ (.A(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\fifo0.fifo_store[33][0] ),
    .A1(_05721_),
    .S(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_05724_),
    .X(_01479_));
 sky130_fd_sc_hd__clkbuf_4 _10866_ (.A(_03872_),
    .X(_05725_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\fifo0.fifo_store[33][1] ),
    .A1(_05725_),
    .S(_05723_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _10868_ (.A(_05726_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(\fifo0.fifo_store[33][2] ),
    .A1(_05493_),
    .S(_05723_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _10870_ (.A(_05727_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(\fifo0.fifo_store[33][3] ),
    .A1(_05495_),
    .S(_05723_),
    .X(_05728_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(_05728_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(\fifo0.fifo_store[33][4] ),
    .A1(_05497_),
    .S(_05723_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _10874_ (.A(_05729_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(\fifo0.fifo_store[33][5] ),
    .A1(_05652_),
    .S(_05723_),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _10876_ (.A(_05730_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(\fifo0.fifo_store[33][6] ),
    .A1(_05500_),
    .S(_05723_),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_1 _10878_ (.A(_05731_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(\fifo0.fifo_store[33][7] ),
    .A1(_05655_),
    .S(_05723_),
    .X(_05732_));
 sky130_fd_sc_hd__clkbuf_1 _10880_ (.A(_05732_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(\fifo0.fifo_store[33][8] ),
    .A1(_05503_),
    .S(_05723_),
    .X(_05733_));
 sky130_fd_sc_hd__clkbuf_1 _10882_ (.A(_05733_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(\fifo0.fifo_store[33][9] ),
    .A1(_05505_),
    .S(_05723_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(_05734_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\fifo0.fifo_store[33][10] ),
    .A1(_05659_),
    .S(_05722_),
    .X(_05735_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_05735_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\fifo0.fifo_store[33][11] ),
    .A1(_05661_),
    .S(_05722_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_05736_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\fifo0.fifo_store[33][12] ),
    .A1(_05509_),
    .S(_05722_),
    .X(_05737_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_05737_),
    .X(_01491_));
 sky130_fd_sc_hd__buf_6 _10891_ (.A(_03908_),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(\fifo0.fifo_store[33][13] ),
    .A1(_05738_),
    .S(_05722_),
    .X(_05739_));
 sky130_fd_sc_hd__clkbuf_1 _10893_ (.A(_05739_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(\fifo0.fifo_store[33][14] ),
    .A1(_05512_),
    .S(_05722_),
    .X(_05740_));
 sky130_fd_sc_hd__clkbuf_1 _10895_ (.A(_05740_),
    .X(_01493_));
 sky130_fd_sc_hd__buf_4 _10896_ (.A(_03914_),
    .X(_05741_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\fifo0.fifo_store[33][15] ),
    .A1(_05741_),
    .S(_05722_),
    .X(_05742_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_05742_),
    .X(_01494_));
 sky130_fd_sc_hd__nor2_8 _10899_ (.A(_04031_),
    .B(_04172_),
    .Y(_05743_));
 sky130_fd_sc_hd__buf_12 _10900_ (.A(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\fifo0.fifo_store[89][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_05745_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\fifo0.fifo_store[89][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_05744_),
    .X(_05746_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_05746_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\fifo0.fifo_store[89][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_05744_),
    .X(_05747_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_05747_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\fifo0.fifo_store[89][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_05744_),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_05748_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\fifo0.fifo_store[89][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_05744_),
    .X(_05749_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_05749_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\fifo0.fifo_store[89][5] ),
    .A1(_05652_),
    .S(_05744_),
    .X(_05750_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_05750_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(\fifo0.fifo_store[89][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_05744_),
    .X(_05751_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_05751_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(\fifo0.fifo_store[89][7] ),
    .A1(_05655_),
    .S(_05744_),
    .X(_05752_));
 sky130_fd_sc_hd__clkbuf_1 _10916_ (.A(_05752_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(\fifo0.fifo_store[89][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_05744_),
    .X(_05753_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(_05753_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(\fifo0.fifo_store[89][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_05744_),
    .X(_05754_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(_05754_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(\fifo0.fifo_store[89][10] ),
    .A1(_05659_),
    .S(_05743_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_1 _10922_ (.A(_05755_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(\fifo0.fifo_store[89][11] ),
    .A1(_05661_),
    .S(_05743_),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_1 _10924_ (.A(_05756_),
    .X(_01506_));
 sky130_fd_sc_hd__buf_4 _10925_ (.A(_03905_),
    .X(_05757_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\fifo0.fifo_store[89][12] ),
    .A1(_05757_),
    .S(_05743_),
    .X(_05758_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_05758_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\fifo0.fifo_store[89][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_05743_),
    .X(_05759_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_05759_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\fifo0.fifo_store[89][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_05743_),
    .X(_05760_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_05760_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\fifo0.fifo_store[89][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_05743_),
    .X(_05761_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(_05761_),
    .X(_01510_));
 sky130_fd_sc_hd__nor2_4 _10934_ (.A(_03815_),
    .B(_05588_),
    .Y(_05762_));
 sky130_fd_sc_hd__buf_6 _10935_ (.A(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\fifo0.fifo_store[32][0] ),
    .A1(_05721_),
    .S(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_1 _10937_ (.A(_05764_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(\fifo0.fifo_store[32][1] ),
    .A1(_05725_),
    .S(_05763_),
    .X(_05765_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(_05765_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_4 _10940_ (.A(_03875_),
    .X(_05766_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\fifo0.fifo_store[32][2] ),
    .A1(_05766_),
    .S(_05763_),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_05767_),
    .X(_01513_));
 sky130_fd_sc_hd__clkbuf_4 _10943_ (.A(_03878_),
    .X(_05768_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(\fifo0.fifo_store[32][3] ),
    .A1(_05768_),
    .S(_05763_),
    .X(_05769_));
 sky130_fd_sc_hd__clkbuf_1 _10945_ (.A(_05769_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_4 _10946_ (.A(_03881_),
    .X(_05770_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\fifo0.fifo_store[32][4] ),
    .A1(_05770_),
    .S(_05763_),
    .X(_05771_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_05771_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\fifo0.fifo_store[32][5] ),
    .A1(_05652_),
    .S(_05763_),
    .X(_05772_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_05772_),
    .X(_01516_));
 sky130_fd_sc_hd__buf_4 _10951_ (.A(_03887_),
    .X(_05773_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(\fifo0.fifo_store[32][6] ),
    .A1(_05773_),
    .S(_05763_),
    .X(_05774_));
 sky130_fd_sc_hd__clkbuf_1 _10953_ (.A(_05774_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10954_ (.A0(\fifo0.fifo_store[32][7] ),
    .A1(_05655_),
    .S(_05763_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _10955_ (.A(_05775_),
    .X(_01518_));
 sky130_fd_sc_hd__buf_4 _10956_ (.A(_03893_),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\fifo0.fifo_store[32][8] ),
    .A1(_05776_),
    .S(_05763_),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_05777_),
    .X(_01519_));
 sky130_fd_sc_hd__clkbuf_4 _10959_ (.A(_03896_),
    .X(_05778_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(\fifo0.fifo_store[32][9] ),
    .A1(_05778_),
    .S(_05763_),
    .X(_05779_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(_05779_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\fifo0.fifo_store[32][10] ),
    .A1(_05659_),
    .S(_05762_),
    .X(_05780_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_05780_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\fifo0.fifo_store[32][11] ),
    .A1(_05661_),
    .S(_05762_),
    .X(_05781_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_05781_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\fifo0.fifo_store[32][12] ),
    .A1(_05757_),
    .S(_05762_),
    .X(_05782_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_05782_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\fifo0.fifo_store[32][13] ),
    .A1(_05738_),
    .S(_05762_),
    .X(_05783_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_05783_),
    .X(_01524_));
 sky130_fd_sc_hd__buf_6 _10970_ (.A(_03911_),
    .X(_05784_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(\fifo0.fifo_store[32][14] ),
    .A1(_05784_),
    .S(_05762_),
    .X(_05785_));
 sky130_fd_sc_hd__clkbuf_1 _10972_ (.A(_05785_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(\fifo0.fifo_store[32][15] ),
    .A1(_05741_),
    .S(_05762_),
    .X(_05786_));
 sky130_fd_sc_hd__clkbuf_1 _10974_ (.A(_05786_),
    .X(_01526_));
 sky130_fd_sc_hd__or2_1 _10975_ (.A(_03812_),
    .B(_04170_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_12 _10976_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__nor2_8 _10977_ (.A(_03920_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__buf_8 _10978_ (.A(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\fifo0.fifo_store[31][0] ),
    .A1(_05721_),
    .S(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(_05791_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\fifo0.fifo_store[31][1] ),
    .A1(_05725_),
    .S(_05790_),
    .X(_05792_));
 sky130_fd_sc_hd__clkbuf_1 _10982_ (.A(_05792_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\fifo0.fifo_store[31][2] ),
    .A1(_05766_),
    .S(_05790_),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_1 _10984_ (.A(_05793_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(\fifo0.fifo_store[31][3] ),
    .A1(_05768_),
    .S(_05790_),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _10986_ (.A(_05794_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\fifo0.fifo_store[31][4] ),
    .A1(_05770_),
    .S(_05790_),
    .X(_05795_));
 sky130_fd_sc_hd__clkbuf_1 _10988_ (.A(_05795_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(\fifo0.fifo_store[31][5] ),
    .A1(_05652_),
    .S(_05790_),
    .X(_05796_));
 sky130_fd_sc_hd__clkbuf_1 _10990_ (.A(_05796_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\fifo0.fifo_store[31][6] ),
    .A1(_05773_),
    .S(_05790_),
    .X(_05797_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_05797_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\fifo0.fifo_store[31][7] ),
    .A1(_05655_),
    .S(_05790_),
    .X(_05798_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(_05798_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\fifo0.fifo_store[31][8] ),
    .A1(_05776_),
    .S(_05790_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(_05799_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\fifo0.fifo_store[31][9] ),
    .A1(_05778_),
    .S(_05790_),
    .X(_05800_));
 sky130_fd_sc_hd__clkbuf_1 _10998_ (.A(_05800_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\fifo0.fifo_store[31][10] ),
    .A1(_05659_),
    .S(_05789_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _11000_ (.A(_05801_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\fifo0.fifo_store[31][11] ),
    .A1(_05661_),
    .S(_05789_),
    .X(_05802_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(_05802_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\fifo0.fifo_store[31][12] ),
    .A1(_05757_),
    .S(_05789_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_05803_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\fifo0.fifo_store[31][13] ),
    .A1(_05738_),
    .S(_05789_),
    .X(_05804_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_05804_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\fifo0.fifo_store[31][14] ),
    .A1(_05784_),
    .S(_05789_),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_05805_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\fifo0.fifo_store[31][15] ),
    .A1(_05741_),
    .S(_05789_),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_05806_),
    .X(_01542_));
 sky130_fd_sc_hd__or2_1 _11011_ (.A(_03943_),
    .B(_05788_),
    .X(_05807_));
 sky130_fd_sc_hd__buf_4 _11012_ (.A(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__buf_8 _11013_ (.A(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[30][0] ),
    .S(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__clkbuf_1 _11015_ (.A(_05810_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[30][1] ),
    .S(_05809_),
    .X(_05811_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(_05811_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[30][2] ),
    .S(_05809_),
    .X(_05812_));
 sky130_fd_sc_hd__clkbuf_1 _11019_ (.A(_05812_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[30][3] ),
    .S(_05809_),
    .X(_05813_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_05813_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[30][4] ),
    .S(_05809_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_1 _11023_ (.A(_05814_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[30][5] ),
    .S(_05809_),
    .X(_05815_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_05815_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[30][6] ),
    .S(_05809_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _11027_ (.A(_05816_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[30][7] ),
    .S(_05809_),
    .X(_05817_));
 sky130_fd_sc_hd__clkbuf_1 _11029_ (.A(_05817_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[30][8] ),
    .S(_05809_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_1 _11031_ (.A(_05818_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[30][9] ),
    .S(_05809_),
    .X(_05819_));
 sky130_fd_sc_hd__clkbuf_1 _11033_ (.A(_05819_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[30][10] ),
    .S(_05808_),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_1 _11035_ (.A(_05820_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[30][11] ),
    .S(_05808_),
    .X(_05821_));
 sky130_fd_sc_hd__clkbuf_1 _11037_ (.A(_05821_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[30][12] ),
    .S(_05808_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_1 _11039_ (.A(_05822_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[30][13] ),
    .S(_05808_),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_1 _11041_ (.A(_05823_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[30][14] ),
    .S(_05808_),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _11043_ (.A(_05824_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[30][15] ),
    .S(_05808_),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_1 _11045_ (.A(_05825_),
    .X(_01558_));
 sky130_fd_sc_hd__nor2_8 _11046_ (.A(_04010_),
    .B(_05788_),
    .Y(_05826_));
 sky130_fd_sc_hd__buf_8 _11047_ (.A(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__mux2_1 _11048_ (.A0(\fifo0.fifo_store[28][0] ),
    .A1(_05721_),
    .S(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_1 _11049_ (.A(_05828_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(\fifo0.fifo_store[28][1] ),
    .A1(_05725_),
    .S(_05827_),
    .X(_05829_));
 sky130_fd_sc_hd__clkbuf_1 _11051_ (.A(_05829_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(\fifo0.fifo_store[28][2] ),
    .A1(_05766_),
    .S(_05827_),
    .X(_05830_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(_05830_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(\fifo0.fifo_store[28][3] ),
    .A1(_05768_),
    .S(_05827_),
    .X(_05831_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_05831_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\fifo0.fifo_store[28][4] ),
    .A1(_05770_),
    .S(_05827_),
    .X(_05832_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(_05832_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\fifo0.fifo_store[28][5] ),
    .A1(_05652_),
    .S(_05827_),
    .X(_05833_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(_05833_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(\fifo0.fifo_store[28][6] ),
    .A1(_05773_),
    .S(_05827_),
    .X(_05834_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_05834_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\fifo0.fifo_store[28][7] ),
    .A1(_05655_),
    .S(_05827_),
    .X(_05835_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_05835_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\fifo0.fifo_store[28][8] ),
    .A1(_05776_),
    .S(_05827_),
    .X(_05836_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_05836_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\fifo0.fifo_store[28][9] ),
    .A1(_05778_),
    .S(_05827_),
    .X(_05837_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_05837_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\fifo0.fifo_store[28][10] ),
    .A1(_05659_),
    .S(_05826_),
    .X(_05838_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_05838_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\fifo0.fifo_store[28][11] ),
    .A1(_05661_),
    .S(_05826_),
    .X(_05839_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(_05839_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(\fifo0.fifo_store[28][12] ),
    .A1(_05757_),
    .S(_05826_),
    .X(_05840_));
 sky130_fd_sc_hd__clkbuf_1 _11073_ (.A(_05840_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(\fifo0.fifo_store[28][13] ),
    .A1(_05738_),
    .S(_05826_),
    .X(_05841_));
 sky130_fd_sc_hd__clkbuf_1 _11075_ (.A(_05841_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(\fifo0.fifo_store[28][14] ),
    .A1(_05784_),
    .S(_05826_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_1 _11077_ (.A(_05842_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(\fifo0.fifo_store[28][15] ),
    .A1(_05741_),
    .S(_05826_),
    .X(_05843_));
 sky130_fd_sc_hd__clkbuf_1 _11079_ (.A(_05843_),
    .X(_01574_));
 sky130_fd_sc_hd__nor2_8 _11080_ (.A(_03814_),
    .B(_03990_),
    .Y(_05844_));
 sky130_fd_sc_hd__buf_6 _11081_ (.A(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(\fifo0.fifo_store[2][0] ),
    .A1(_05721_),
    .S(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__clkbuf_1 _11083_ (.A(_05846_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(\fifo0.fifo_store[2][1] ),
    .A1(_05725_),
    .S(_05845_),
    .X(_05847_));
 sky130_fd_sc_hd__clkbuf_1 _11085_ (.A(_05847_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(\fifo0.fifo_store[2][2] ),
    .A1(_05766_),
    .S(_05845_),
    .X(_05848_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(_05848_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(\fifo0.fifo_store[2][3] ),
    .A1(_05768_),
    .S(_05845_),
    .X(_05849_));
 sky130_fd_sc_hd__clkbuf_1 _11089_ (.A(_05849_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(\fifo0.fifo_store[2][4] ),
    .A1(_05770_),
    .S(_05845_),
    .X(_05850_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(_05850_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\fifo0.fifo_store[2][5] ),
    .A1(_05652_),
    .S(_05845_),
    .X(_05851_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_05851_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\fifo0.fifo_store[2][6] ),
    .A1(_05773_),
    .S(_05845_),
    .X(_05852_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_05852_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\fifo0.fifo_store[2][7] ),
    .A1(_05655_),
    .S(_05845_),
    .X(_05853_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_05853_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\fifo0.fifo_store[2][8] ),
    .A1(_05776_),
    .S(_05845_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_05854_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\fifo0.fifo_store[2][9] ),
    .A1(_05778_),
    .S(_05845_),
    .X(_05855_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_05855_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(\fifo0.fifo_store[2][10] ),
    .A1(_05659_),
    .S(_05844_),
    .X(_05856_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(_05856_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(\fifo0.fifo_store[2][11] ),
    .A1(_05661_),
    .S(_05844_),
    .X(_05857_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(_05857_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(\fifo0.fifo_store[2][12] ),
    .A1(_05757_),
    .S(_05844_),
    .X(_05858_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(_05858_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\fifo0.fifo_store[2][13] ),
    .A1(_05738_),
    .S(_05844_),
    .X(_05859_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(_05859_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(\fifo0.fifo_store[2][14] ),
    .A1(_05784_),
    .S(_05844_),
    .X(_05860_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_05860_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(\fifo0.fifo_store[2][15] ),
    .A1(_05741_),
    .S(_05844_),
    .X(_05861_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(_05861_),
    .X(_01590_));
 sky130_fd_sc_hd__nor2_8 _11114_ (.A(_03920_),
    .B(_04356_),
    .Y(_05862_));
 sky130_fd_sc_hd__buf_8 _11115_ (.A(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(\fifo0.fifo_store[15][0] ),
    .A1(_05721_),
    .S(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__clkbuf_1 _11117_ (.A(_05864_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(\fifo0.fifo_store[15][1] ),
    .A1(_05725_),
    .S(_05863_),
    .X(_05865_));
 sky130_fd_sc_hd__clkbuf_1 _11119_ (.A(_05865_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(\fifo0.fifo_store[15][2] ),
    .A1(_05766_),
    .S(_05863_),
    .X(_05866_));
 sky130_fd_sc_hd__clkbuf_1 _11121_ (.A(_05866_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _11122_ (.A0(\fifo0.fifo_store[15][3] ),
    .A1(_05768_),
    .S(_05863_),
    .X(_05867_));
 sky130_fd_sc_hd__clkbuf_1 _11123_ (.A(_05867_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\fifo0.fifo_store[15][4] ),
    .A1(_05770_),
    .S(_05863_),
    .X(_05868_));
 sky130_fd_sc_hd__clkbuf_1 _11125_ (.A(_05868_),
    .X(_01595_));
 sky130_fd_sc_hd__buf_4 _11126_ (.A(_03838_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(\fifo0.fifo_store[15][5] ),
    .A1(_05869_),
    .S(_05863_),
    .X(_05870_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(_05870_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(\fifo0.fifo_store[15][6] ),
    .A1(_05773_),
    .S(_05863_),
    .X(_05871_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_05871_),
    .X(_01597_));
 sky130_fd_sc_hd__buf_4 _11131_ (.A(_03843_),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(\fifo0.fifo_store[15][7] ),
    .A1(_05872_),
    .S(_05863_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _11133_ (.A(_05873_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(\fifo0.fifo_store[15][8] ),
    .A1(_05776_),
    .S(_05863_),
    .X(_05874_));
 sky130_fd_sc_hd__clkbuf_1 _11135_ (.A(_05874_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(\fifo0.fifo_store[15][9] ),
    .A1(_05778_),
    .S(_05863_),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(_05875_),
    .X(_01600_));
 sky130_fd_sc_hd__clkbuf_4 _11138_ (.A(_03850_),
    .X(_05876_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(\fifo0.fifo_store[15][10] ),
    .A1(_05876_),
    .S(_05862_),
    .X(_05877_));
 sky130_fd_sc_hd__clkbuf_1 _11140_ (.A(_05877_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_4 _11141_ (.A(_03853_),
    .X(_05878_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(\fifo0.fifo_store[15][11] ),
    .A1(_05878_),
    .S(_05862_),
    .X(_05879_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_05879_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(\fifo0.fifo_store[15][12] ),
    .A1(_05757_),
    .S(_05862_),
    .X(_05880_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(_05880_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(\fifo0.fifo_store[15][13] ),
    .A1(_05738_),
    .S(_05862_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(_05881_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(\fifo0.fifo_store[15][14] ),
    .A1(_05784_),
    .S(_05862_),
    .X(_05882_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(_05882_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(\fifo0.fifo_store[15][15] ),
    .A1(_05741_),
    .S(_05862_),
    .X(_05883_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(_05883_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_4 _11152_ (.A(_03814_),
    .B(_04277_),
    .Y(_05884_));
 sky130_fd_sc_hd__buf_6 _11153_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(\fifo0.fifo_store[4][0] ),
    .A1(_05721_),
    .S(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_05886_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(\fifo0.fifo_store[4][1] ),
    .A1(_05725_),
    .S(_05885_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_1 _11157_ (.A(_05887_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(\fifo0.fifo_store[4][2] ),
    .A1(_05766_),
    .S(_05885_),
    .X(_05888_));
 sky130_fd_sc_hd__clkbuf_1 _11159_ (.A(_05888_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(\fifo0.fifo_store[4][3] ),
    .A1(_05768_),
    .S(_05885_),
    .X(_05889_));
 sky130_fd_sc_hd__clkbuf_1 _11161_ (.A(_05889_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(\fifo0.fifo_store[4][4] ),
    .A1(_05770_),
    .S(_05885_),
    .X(_05890_));
 sky130_fd_sc_hd__clkbuf_1 _11163_ (.A(_05890_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _11164_ (.A0(\fifo0.fifo_store[4][5] ),
    .A1(_05869_),
    .S(_05885_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_1 _11165_ (.A(_05891_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(\fifo0.fifo_store[4][6] ),
    .A1(_05773_),
    .S(_05885_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_1 _11167_ (.A(_05892_),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _11168_ (.A0(\fifo0.fifo_store[4][7] ),
    .A1(_05872_),
    .S(_05885_),
    .X(_05893_));
 sky130_fd_sc_hd__clkbuf_1 _11169_ (.A(_05893_),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _11170_ (.A0(\fifo0.fifo_store[4][8] ),
    .A1(_05776_),
    .S(_05885_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _11171_ (.A(_05894_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(\fifo0.fifo_store[4][9] ),
    .A1(_05778_),
    .S(_05885_),
    .X(_05895_));
 sky130_fd_sc_hd__clkbuf_1 _11173_ (.A(_05895_),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(\fifo0.fifo_store[4][10] ),
    .A1(_05876_),
    .S(_05884_),
    .X(_05896_));
 sky130_fd_sc_hd__clkbuf_1 _11175_ (.A(_05896_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _11176_ (.A0(\fifo0.fifo_store[4][11] ),
    .A1(_05878_),
    .S(_05884_),
    .X(_05897_));
 sky130_fd_sc_hd__clkbuf_1 _11177_ (.A(_05897_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(\fifo0.fifo_store[4][12] ),
    .A1(_05757_),
    .S(_05884_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(_05898_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(\fifo0.fifo_store[4][13] ),
    .A1(_05738_),
    .S(_05884_),
    .X(_05899_));
 sky130_fd_sc_hd__clkbuf_1 _11181_ (.A(_05899_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(\fifo0.fifo_store[4][14] ),
    .A1(_05784_),
    .S(_05884_),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_1 _11183_ (.A(_05900_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(\fifo0.fifo_store[4][15] ),
    .A1(_05741_),
    .S(_05884_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_05901_),
    .X(_01622_));
 sky130_fd_sc_hd__buf_4 _11186_ (.A(net21),
    .X(_05902_));
 sky130_fd_sc_hd__buf_4 _11187_ (.A(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__and2_1 _11188_ (.A(_05903_),
    .B(net1),
    .X(_05904_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_05904_),
    .X(_01623_));
 sky130_fd_sc_hd__clkbuf_4 _11190_ (.A(net21),
    .X(_05905_));
 sky130_fd_sc_hd__and2_1 _11191_ (.A(_05905_),
    .B(net8),
    .X(_05906_));
 sky130_fd_sc_hd__clkbuf_1 _11192_ (.A(_05906_),
    .X(_01624_));
 sky130_fd_sc_hd__and2_1 _11193_ (.A(_05905_),
    .B(net9),
    .X(_05907_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_05907_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_1 _11195_ (.A(_05905_),
    .B(net10),
    .X(_05908_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(_05908_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_1 _11197_ (.A(_05905_),
    .B(net11),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_1 _11198_ (.A(_05909_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_1 _11199_ (.A(_05905_),
    .B(net12),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(_05910_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_1 _11201_ (.A(_05905_),
    .B(net13),
    .X(_05911_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(_05911_),
    .X(_01629_));
 sky130_fd_sc_hd__and2_1 _11203_ (.A(_05905_),
    .B(net14),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(_05912_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_1 _11205_ (.A(_05905_),
    .B(net15),
    .X(_05913_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(_05913_),
    .X(_01631_));
 sky130_fd_sc_hd__and2_1 _11207_ (.A(_05905_),
    .B(net16),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_05914_),
    .X(_01632_));
 sky130_fd_sc_hd__and2_1 _11209_ (.A(_05905_),
    .B(net2),
    .X(_05915_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_05915_),
    .X(_01633_));
 sky130_fd_sc_hd__buf_4 _11211_ (.A(net21),
    .X(_05916_));
 sky130_fd_sc_hd__and2_1 _11212_ (.A(_05916_),
    .B(net3),
    .X(_05917_));
 sky130_fd_sc_hd__clkbuf_1 _11213_ (.A(_05917_),
    .X(_01634_));
 sky130_fd_sc_hd__and2_1 _11214_ (.A(_05916_),
    .B(net4),
    .X(_05918_));
 sky130_fd_sc_hd__clkbuf_1 _11215_ (.A(_05918_),
    .X(_01635_));
 sky130_fd_sc_hd__and2_1 _11216_ (.A(_05916_),
    .B(net5),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _11217_ (.A(_05919_),
    .X(_01636_));
 sky130_fd_sc_hd__and2_1 _11218_ (.A(_05916_),
    .B(net6),
    .X(_05920_));
 sky130_fd_sc_hd__clkbuf_1 _11219_ (.A(_05920_),
    .X(_01637_));
 sky130_fd_sc_hd__and2_1 _11220_ (.A(_05916_),
    .B(net7),
    .X(_05921_));
 sky130_fd_sc_hd__clkbuf_1 _11221_ (.A(_05921_),
    .X(_01638_));
 sky130_fd_sc_hd__and2_1 _11222_ (.A(_05916_),
    .B(\fifo0.fifo_rdy_del1 ),
    .X(_05922_));
 sky130_fd_sc_hd__clkbuf_1 _11223_ (.A(_05922_),
    .X(_01639_));
 sky130_fd_sc_hd__and2_1 _11224_ (.A(_05916_),
    .B(net17),
    .X(_05923_));
 sky130_fd_sc_hd__clkbuf_1 _11225_ (.A(_05923_),
    .X(_01640_));
 sky130_fd_sc_hd__buf_4 _11226_ (.A(_03799_),
    .X(_05924_));
 sky130_fd_sc_hd__nor2_1 _11227_ (.A(_05924_),
    .B(\dsmod0.fetch_ctr[0] ),
    .Y(_01641_));
 sky130_fd_sc_hd__nor2_1 _11228_ (.A(\dsmod0.fetch_ctr[1] ),
    .B(\dsmod0.fetch_ctr[0] ),
    .Y(_05925_));
 sky130_fd_sc_hd__and2_1 _11229_ (.A(\dsmod0.fetch_ctr[1] ),
    .B(\dsmod0.fetch_ctr[0] ),
    .X(_05926_));
 sky130_fd_sc_hd__buf_4 _11230_ (.A(_05902_),
    .X(_05927_));
 sky130_fd_sc_hd__o21a_1 _11231_ (.A1(_05925_),
    .A2(_05926_),
    .B1(_05927_),
    .X(_01642_));
 sky130_fd_sc_hd__and2b_1 _11232_ (.A_N(\dsmod0.fetch_ctr[2] ),
    .B(_05925_),
    .X(_05928_));
 sky130_fd_sc_hd__o21a_1 _11233_ (.A1(\dsmod0.fetch_ctr[1] ),
    .A2(\dsmod0.fetch_ctr[0] ),
    .B1(\dsmod0.fetch_ctr[2] ),
    .X(_05929_));
 sky130_fd_sc_hd__o21a_1 _11234_ (.A1(_05928_),
    .A2(_05929_),
    .B1(_05927_),
    .X(_01643_));
 sky130_fd_sc_hd__or4_2 _11235_ (.A(\dsmod0.fetch_ctr[1] ),
    .B(\dsmod0.fetch_ctr[0] ),
    .C(\dsmod0.fetch_ctr[3] ),
    .D(\dsmod0.fetch_ctr[2] ),
    .X(_05930_));
 sky130_fd_sc_hd__or2b_1 _11236_ (.A(_05928_),
    .B_N(\dsmod0.fetch_ctr[3] ),
    .X(_05931_));
 sky130_fd_sc_hd__a21oi_1 _11237_ (.A1(_05930_),
    .A2(_05931_),
    .B1(_05924_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _11238_ (.A(\dsmod0.fetch_ctr[4] ),
    .B(_05930_),
    .Y(_05932_));
 sky130_fd_sc_hd__and2_1 _11239_ (.A(\dsmod0.fetch_ctr[4] ),
    .B(_05930_),
    .X(_05933_));
 sky130_fd_sc_hd__o21a_1 _11240_ (.A1(_05932_),
    .A2(_05933_),
    .B1(_05927_),
    .X(_01645_));
 sky130_fd_sc_hd__or4_1 _11241_ (.A(\dsmod0.fetch_ctr[5] ),
    .B(\dsmod0.fetch_ctr[4] ),
    .C(\dsmod0.fetch_ctr[6] ),
    .D(_05930_),
    .X(_05934_));
 sky130_fd_sc_hd__nor2_2 _11242_ (.A(\dsmod0.fetch_ctr[7] ),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__inv_2 _11243_ (.A(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__xor2_1 _11244_ (.A(\dsmod0.fetch_ctr[5] ),
    .B(_05932_),
    .X(_05937_));
 sky130_fd_sc_hd__o311a_1 _11245_ (.A1(net19),
    .A2(net20),
    .A3(_05936_),
    .B1(_05937_),
    .C1(_05903_),
    .X(_01646_));
 sky130_fd_sc_hd__o31a_1 _11246_ (.A1(\dsmod0.fetch_ctr[5] ),
    .A2(\dsmod0.fetch_ctr[4] ),
    .A3(_05930_),
    .B1(\dsmod0.fetch_ctr[6] ),
    .X(_05938_));
 sky130_fd_sc_hd__o21ba_1 _11247_ (.A1(\dsmod0.fetch_ctr[7] ),
    .A2(net20),
    .B1_N(_05934_),
    .X(_05939_));
 sky130_fd_sc_hd__o21a_1 _11248_ (.A1(_05938_),
    .A2(_05939_),
    .B1(_05927_),
    .X(_01647_));
 sky130_fd_sc_hd__and3_1 _11249_ (.A(net19),
    .B(net20),
    .C(_05935_),
    .X(_05940_));
 sky130_fd_sc_hd__a21oi_1 _11250_ (.A1(\dsmod0.fetch_ctr[7] ),
    .A2(_05934_),
    .B1(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(_05924_),
    .B(_05941_),
    .Y(_01648_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(_03819_),
    .A1(_03824_),
    .S(\fifo0.write_ptr[0] ),
    .X(_05942_));
 sky130_fd_sc_hd__clkbuf_1 _11253_ (.A(_05942_),
    .X(_01649_));
 sky130_fd_sc_hd__a21bo_1 _11254_ (.A1(\fifo0.write_ptr[1] ),
    .A2(_03824_),
    .B1_N(_03917_),
    .X(_01650_));
 sky130_fd_sc_hd__a21bo_1 _11255_ (.A1(\fifo0.write_ptr[2] ),
    .A2(_03824_),
    .B1_N(_03942_),
    .X(_01651_));
 sky130_fd_sc_hd__a21o_1 _11256_ (.A1(\fifo0.write_ptr[3] ),
    .A2(_03824_),
    .B1(_03804_),
    .X(_01652_));
 sky130_fd_sc_hd__a21o_1 _11257_ (.A1(\fifo0.write_ptr[4] ),
    .A2(_03824_),
    .B1(_03805_),
    .X(_01653_));
 sky130_fd_sc_hd__a21o_1 _11258_ (.A1(\fifo0.write_ptr[5] ),
    .A2(_03824_),
    .B1(_03809_),
    .X(_01654_));
 sky130_fd_sc_hd__a21o_1 _11259_ (.A1(\fifo0.write_ptr[6] ),
    .A2(_03824_),
    .B1(_03811_),
    .X(_01655_));
 sky130_fd_sc_hd__o21a_2 _11260_ (.A1(net22),
    .A2(_03779_),
    .B1(_05935_),
    .X(_05943_));
 sky130_fd_sc_hd__and2_1 _11261_ (.A(\fifo0.read_ptr[0] ),
    .B(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__o21ai_1 _11262_ (.A1(\fifo0.read_ptr[0] ),
    .A2(_05943_),
    .B1(_05903_),
    .Y(_05945_));
 sky130_fd_sc_hd__nor2_1 _11263_ (.A(_05944_),
    .B(_05945_),
    .Y(_01656_));
 sky130_fd_sc_hd__and3_1 _11264_ (.A(\fifo0.read_ptr[1] ),
    .B(\fifo0.read_ptr[0] ),
    .C(_05943_),
    .X(_05946_));
 sky130_fd_sc_hd__o21ai_1 _11265_ (.A1(\fifo0.read_ptr[1] ),
    .A2(_05944_),
    .B1(_05903_),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _11266_ (.A(_05946_),
    .B(_05947_),
    .Y(_01657_));
 sky130_fd_sc_hd__and3_1 _11267_ (.A(\fifo0.read_ptr[2] ),
    .B(\fifo0.read_ptr[1] ),
    .C(_05944_),
    .X(_05948_));
 sky130_fd_sc_hd__o21ai_1 _11268_ (.A1(\fifo0.read_ptr[2] ),
    .A2(_05946_),
    .B1(_05903_),
    .Y(_05949_));
 sky130_fd_sc_hd__nor2_1 _11269_ (.A(_05948_),
    .B(_05949_),
    .Y(_01658_));
 sky130_fd_sc_hd__and2_1 _11270_ (.A(\fifo0.read_ptr[3] ),
    .B(_05948_),
    .X(_05950_));
 sky130_fd_sc_hd__o21ai_1 _11271_ (.A1(\fifo0.read_ptr[3] ),
    .A2(_05948_),
    .B1(_05903_),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2_1 _11272_ (.A(_05950_),
    .B(_05951_),
    .Y(_01659_));
 sky130_fd_sc_hd__and3_1 _11273_ (.A(\fifo0.read_ptr[4] ),
    .B(\fifo0.read_ptr[3] ),
    .C(_05948_),
    .X(_05952_));
 sky130_fd_sc_hd__o21ai_1 _11274_ (.A1(\fifo0.read_ptr[4] ),
    .A2(_05950_),
    .B1(_05903_),
    .Y(_05953_));
 sky130_fd_sc_hd__nor2_1 _11275_ (.A(_05952_),
    .B(_05953_),
    .Y(_01660_));
 sky130_fd_sc_hd__and2_1 _11276_ (.A(\fifo0.read_ptr[5] ),
    .B(_05952_),
    .X(_05954_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11277_ (.A(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__o21ai_1 _11278_ (.A1(\fifo0.read_ptr[5] ),
    .A2(_05952_),
    .B1(_05903_),
    .Y(_05956_));
 sky130_fd_sc_hd__nor2_1 _11279_ (.A(_05955_),
    .B(_05956_),
    .Y(_01661_));
 sky130_fd_sc_hd__o21ai_1 _11280_ (.A1(\fifo0.read_ptr[6] ),
    .A2(_05955_),
    .B1(_05903_),
    .Y(_05957_));
 sky130_fd_sc_hd__a21oi_1 _11281_ (.A1(\fifo0.read_ptr[6] ),
    .A2(_05955_),
    .B1(_05957_),
    .Y(_01662_));
 sky130_fd_sc_hd__o211a_1 _11282_ (.A1(net36),
    .A2(_03798_),
    .B1(_05903_),
    .C1(\fifo0.fifo_rdy ),
    .X(_01663_));
 sky130_fd_sc_hd__nor2_8 _11283_ (.A(_04052_),
    .B(_05001_),
    .Y(_05958_));
 sky130_fd_sc_hd__buf_6 _11284_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(\fifo0.fifo_store[59][0] ),
    .A1(_05721_),
    .S(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__clkbuf_1 _11286_ (.A(_05960_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _11287_ (.A0(\fifo0.fifo_store[59][1] ),
    .A1(_05725_),
    .S(_05959_),
    .X(_05961_));
 sky130_fd_sc_hd__clkbuf_1 _11288_ (.A(_05961_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\fifo0.fifo_store[59][2] ),
    .A1(_05766_),
    .S(_05959_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05962_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(\fifo0.fifo_store[59][3] ),
    .A1(_05768_),
    .S(_05959_),
    .X(_05963_));
 sky130_fd_sc_hd__clkbuf_1 _11292_ (.A(_05963_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(\fifo0.fifo_store[59][4] ),
    .A1(_05770_),
    .S(_05959_),
    .X(_05964_));
 sky130_fd_sc_hd__clkbuf_1 _11294_ (.A(_05964_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(\fifo0.fifo_store[59][5] ),
    .A1(_05869_),
    .S(_05959_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(_05965_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(\fifo0.fifo_store[59][6] ),
    .A1(_05773_),
    .S(_05959_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _11298_ (.A(_05966_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(\fifo0.fifo_store[59][7] ),
    .A1(_05872_),
    .S(_05959_),
    .X(_05967_));
 sky130_fd_sc_hd__clkbuf_1 _11300_ (.A(_05967_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(\fifo0.fifo_store[59][8] ),
    .A1(_05776_),
    .S(_05959_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_05968_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(\fifo0.fifo_store[59][9] ),
    .A1(_05778_),
    .S(_05959_),
    .X(_05969_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(_05969_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(\fifo0.fifo_store[59][10] ),
    .A1(_05876_),
    .S(_05958_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_05970_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(\fifo0.fifo_store[59][11] ),
    .A1(_05878_),
    .S(_05958_),
    .X(_05971_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_05971_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(\fifo0.fifo_store[59][12] ),
    .A1(_05757_),
    .S(_05958_),
    .X(_05972_));
 sky130_fd_sc_hd__clkbuf_1 _11310_ (.A(_05972_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(\fifo0.fifo_store[59][13] ),
    .A1(_05738_),
    .S(_05958_),
    .X(_05973_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_05973_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(\fifo0.fifo_store[59][14] ),
    .A1(_05784_),
    .S(_05958_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_05974_),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(\fifo0.fifo_store[59][15] ),
    .A1(_05741_),
    .S(_05958_),
    .X(_05975_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05975_),
    .X(_01679_));
 sky130_fd_sc_hd__nor2_8 _11317_ (.A(_03964_),
    .B(_04356_),
    .Y(_05976_));
 sky130_fd_sc_hd__buf_8 _11318_ (.A(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(\fifo0.fifo_store[13][0] ),
    .A1(_05721_),
    .S(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__clkbuf_1 _11320_ (.A(_05978_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _11321_ (.A0(\fifo0.fifo_store[13][1] ),
    .A1(_05725_),
    .S(_05977_),
    .X(_05979_));
 sky130_fd_sc_hd__clkbuf_1 _11322_ (.A(_05979_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _11323_ (.A0(\fifo0.fifo_store[13][2] ),
    .A1(_05766_),
    .S(_05977_),
    .X(_05980_));
 sky130_fd_sc_hd__clkbuf_1 _11324_ (.A(_05980_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _11325_ (.A0(\fifo0.fifo_store[13][3] ),
    .A1(_05768_),
    .S(_05977_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_1 _11326_ (.A(_05981_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _11327_ (.A0(\fifo0.fifo_store[13][4] ),
    .A1(_05770_),
    .S(_05977_),
    .X(_05982_));
 sky130_fd_sc_hd__clkbuf_1 _11328_ (.A(_05982_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _11329_ (.A0(\fifo0.fifo_store[13][5] ),
    .A1(_05869_),
    .S(_05977_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _11330_ (.A(_05983_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _11331_ (.A0(\fifo0.fifo_store[13][6] ),
    .A1(_05773_),
    .S(_05977_),
    .X(_05984_));
 sky130_fd_sc_hd__clkbuf_1 _11332_ (.A(_05984_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _11333_ (.A0(\fifo0.fifo_store[13][7] ),
    .A1(_05872_),
    .S(_05977_),
    .X(_05985_));
 sky130_fd_sc_hd__clkbuf_1 _11334_ (.A(_05985_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _11335_ (.A0(\fifo0.fifo_store[13][8] ),
    .A1(_05776_),
    .S(_05977_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _11336_ (.A(_05986_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _11337_ (.A0(\fifo0.fifo_store[13][9] ),
    .A1(_05778_),
    .S(_05977_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _11338_ (.A(_05987_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _11339_ (.A0(\fifo0.fifo_store[13][10] ),
    .A1(_05876_),
    .S(_05976_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _11340_ (.A(_05988_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _11341_ (.A0(\fifo0.fifo_store[13][11] ),
    .A1(_05878_),
    .S(_05976_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _11342_ (.A(_05989_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(\fifo0.fifo_store[13][12] ),
    .A1(_05757_),
    .S(_05976_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_1 _11344_ (.A(_05990_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(\fifo0.fifo_store[13][13] ),
    .A1(_05738_),
    .S(_05976_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _11346_ (.A(_05991_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(\fifo0.fifo_store[13][14] ),
    .A1(_05784_),
    .S(_05976_),
    .X(_05992_));
 sky130_fd_sc_hd__clkbuf_1 _11348_ (.A(_05992_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _11349_ (.A0(\fifo0.fifo_store[13][15] ),
    .A1(_05741_),
    .S(_05976_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _11350_ (.A(_05993_),
    .X(_01695_));
 sky130_fd_sc_hd__or2_1 _11351_ (.A(_03812_),
    .B(_03865_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_12 _11352_ (.A(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__nor2_8 _11353_ (.A(_03815_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__buf_8 _11354_ (.A(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(\fifo0.fifo_store[16][0] ),
    .A1(_05721_),
    .S(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_1 _11356_ (.A(_05998_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _11357_ (.A0(\fifo0.fifo_store[16][1] ),
    .A1(_05725_),
    .S(_05997_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _11358_ (.A(_05999_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _11359_ (.A0(\fifo0.fifo_store[16][2] ),
    .A1(_05766_),
    .S(_05997_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _11360_ (.A(_06000_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(\fifo0.fifo_store[16][3] ),
    .A1(_05768_),
    .S(_05997_),
    .X(_06001_));
 sky130_fd_sc_hd__clkbuf_1 _11362_ (.A(_06001_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _11363_ (.A0(\fifo0.fifo_store[16][4] ),
    .A1(_05770_),
    .S(_05997_),
    .X(_06002_));
 sky130_fd_sc_hd__clkbuf_1 _11364_ (.A(_06002_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(\fifo0.fifo_store[16][5] ),
    .A1(_05869_),
    .S(_05997_),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_1 _11366_ (.A(_06003_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _11367_ (.A0(\fifo0.fifo_store[16][6] ),
    .A1(_05773_),
    .S(_05997_),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_1 _11368_ (.A(_06004_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(\fifo0.fifo_store[16][7] ),
    .A1(_05872_),
    .S(_05997_),
    .X(_06005_));
 sky130_fd_sc_hd__clkbuf_1 _11370_ (.A(_06005_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(\fifo0.fifo_store[16][8] ),
    .A1(_05776_),
    .S(_05997_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _11372_ (.A(_06006_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(\fifo0.fifo_store[16][9] ),
    .A1(_05778_),
    .S(_05997_),
    .X(_06007_));
 sky130_fd_sc_hd__clkbuf_1 _11374_ (.A(_06007_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(\fifo0.fifo_store[16][10] ),
    .A1(_05876_),
    .S(_05996_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_1 _11376_ (.A(_06008_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(\fifo0.fifo_store[16][11] ),
    .A1(_05878_),
    .S(_05996_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_1 _11378_ (.A(_06009_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(\fifo0.fifo_store[16][12] ),
    .A1(_05757_),
    .S(_05996_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_1 _11380_ (.A(_06010_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(\fifo0.fifo_store[16][13] ),
    .A1(_05738_),
    .S(_05996_),
    .X(_06011_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(_06011_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(\fifo0.fifo_store[16][14] ),
    .A1(_05784_),
    .S(_05996_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_1 _11384_ (.A(_06012_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(\fifo0.fifo_store[16][15] ),
    .A1(_05741_),
    .S(_05996_),
    .X(_06013_));
 sky130_fd_sc_hd__clkbuf_1 _11386_ (.A(_06013_),
    .X(_01711_));
 sky130_fd_sc_hd__nor2_8 _11387_ (.A(_04031_),
    .B(_05995_),
    .Y(_06014_));
 sky130_fd_sc_hd__buf_8 _11388_ (.A(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(\fifo0.fifo_store[17][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_1 _11390_ (.A(_06016_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(\fifo0.fifo_store[17][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_06015_),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(_06017_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(\fifo0.fifo_store[17][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_06015_),
    .X(_06018_));
 sky130_fd_sc_hd__clkbuf_1 _11394_ (.A(_06018_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(\fifo0.fifo_store[17][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_06015_),
    .X(_06019_));
 sky130_fd_sc_hd__clkbuf_1 _11396_ (.A(_06019_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _11397_ (.A0(\fifo0.fifo_store[17][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_06015_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _11398_ (.A(_06020_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _11399_ (.A0(\fifo0.fifo_store[17][5] ),
    .A1(_05869_),
    .S(_06015_),
    .X(_06021_));
 sky130_fd_sc_hd__clkbuf_1 _11400_ (.A(_06021_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _11401_ (.A0(\fifo0.fifo_store[17][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_06015_),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_1 _11402_ (.A(_06022_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(\fifo0.fifo_store[17][7] ),
    .A1(_05872_),
    .S(_06015_),
    .X(_06023_));
 sky130_fd_sc_hd__clkbuf_1 _11404_ (.A(_06023_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(\fifo0.fifo_store[17][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_06015_),
    .X(_06024_));
 sky130_fd_sc_hd__clkbuf_1 _11406_ (.A(_06024_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _11407_ (.A0(\fifo0.fifo_store[17][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_06015_),
    .X(_06025_));
 sky130_fd_sc_hd__clkbuf_1 _11408_ (.A(_06025_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _11409_ (.A0(\fifo0.fifo_store[17][10] ),
    .A1(_05876_),
    .S(_06014_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _11410_ (.A(_06026_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _11411_ (.A0(\fifo0.fifo_store[17][11] ),
    .A1(_05878_),
    .S(_06014_),
    .X(_06027_));
 sky130_fd_sc_hd__clkbuf_1 _11412_ (.A(_06027_),
    .X(_01723_));
 sky130_fd_sc_hd__buf_4 _11413_ (.A(_03855_),
    .X(_06028_));
 sky130_fd_sc_hd__mux2_1 _11414_ (.A0(\fifo0.fifo_store[17][12] ),
    .A1(_06028_),
    .S(_06014_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_1 _11415_ (.A(_06029_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(\fifo0.fifo_store[17][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_06014_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_1 _11417_ (.A(_06030_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(\fifo0.fifo_store[17][14] ),
    .A1(\fifo0.fifo_data[14] ),
    .S(_06014_),
    .X(_06031_));
 sky130_fd_sc_hd__clkbuf_1 _11419_ (.A(_06031_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _11420_ (.A0(\fifo0.fifo_store[17][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_06014_),
    .X(_06032_));
 sky130_fd_sc_hd__clkbuf_1 _11421_ (.A(_06032_),
    .X(_01727_));
 sky130_fd_sc_hd__clkbuf_4 _11422_ (.A(_03820_),
    .X(_06033_));
 sky130_fd_sc_hd__nor2_8 _11423_ (.A(_03815_),
    .B(_04690_),
    .Y(_06034_));
 sky130_fd_sc_hd__buf_8 _11424_ (.A(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(\fifo0.fifo_store[48][0] ),
    .A1(_06033_),
    .S(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__clkbuf_1 _11426_ (.A(_06036_),
    .X(_01728_));
 sky130_fd_sc_hd__buf_4 _11427_ (.A(_03872_),
    .X(_06037_));
 sky130_fd_sc_hd__mux2_1 _11428_ (.A0(\fifo0.fifo_store[48][1] ),
    .A1(_06037_),
    .S(_06035_),
    .X(_06038_));
 sky130_fd_sc_hd__clkbuf_1 _11429_ (.A(_06038_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _11430_ (.A0(\fifo0.fifo_store[48][2] ),
    .A1(_05766_),
    .S(_06035_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_1 _11431_ (.A(_06039_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _11432_ (.A0(\fifo0.fifo_store[48][3] ),
    .A1(_05768_),
    .S(_06035_),
    .X(_06040_));
 sky130_fd_sc_hd__clkbuf_1 _11433_ (.A(_06040_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(\fifo0.fifo_store[48][4] ),
    .A1(_05770_),
    .S(_06035_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_1 _11435_ (.A(_06041_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _11436_ (.A0(\fifo0.fifo_store[48][5] ),
    .A1(_05869_),
    .S(_06035_),
    .X(_06042_));
 sky130_fd_sc_hd__clkbuf_1 _11437_ (.A(_06042_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(\fifo0.fifo_store[48][6] ),
    .A1(_05773_),
    .S(_06035_),
    .X(_06043_));
 sky130_fd_sc_hd__clkbuf_1 _11439_ (.A(_06043_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(\fifo0.fifo_store[48][7] ),
    .A1(_05872_),
    .S(_06035_),
    .X(_06044_));
 sky130_fd_sc_hd__clkbuf_1 _11441_ (.A(_06044_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(\fifo0.fifo_store[48][8] ),
    .A1(_05776_),
    .S(_06035_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_06045_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _11444_ (.A0(\fifo0.fifo_store[48][9] ),
    .A1(_05778_),
    .S(_06035_),
    .X(_06046_));
 sky130_fd_sc_hd__clkbuf_1 _11445_ (.A(_06046_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(\fifo0.fifo_store[48][10] ),
    .A1(_05876_),
    .S(_06034_),
    .X(_06047_));
 sky130_fd_sc_hd__clkbuf_1 _11447_ (.A(_06047_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(\fifo0.fifo_store[48][11] ),
    .A1(_05878_),
    .S(_06034_),
    .X(_06048_));
 sky130_fd_sc_hd__clkbuf_1 _11449_ (.A(_06048_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _11450_ (.A0(\fifo0.fifo_store[48][12] ),
    .A1(_06028_),
    .S(_06034_),
    .X(_06049_));
 sky130_fd_sc_hd__clkbuf_1 _11451_ (.A(_06049_),
    .X(_01740_));
 sky130_fd_sc_hd__clkbuf_8 _11452_ (.A(_03908_),
    .X(_06050_));
 sky130_fd_sc_hd__mux2_1 _11453_ (.A0(\fifo0.fifo_store[48][13] ),
    .A1(_06050_),
    .S(_06034_),
    .X(_06051_));
 sky130_fd_sc_hd__clkbuf_1 _11454_ (.A(_06051_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(\fifo0.fifo_store[48][14] ),
    .A1(_05784_),
    .S(_06034_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_1 _11456_ (.A(_06052_),
    .X(_01742_));
 sky130_fd_sc_hd__clkbuf_4 _11457_ (.A(_03914_),
    .X(_06053_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(\fifo0.fifo_store[48][15] ),
    .A1(_06053_),
    .S(_06034_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_1 _11459_ (.A(_06054_),
    .X(_01743_));
 sky130_fd_sc_hd__nor2_8 _11460_ (.A(_04052_),
    .B(_05788_),
    .Y(_06055_));
 sky130_fd_sc_hd__buf_8 _11461_ (.A(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(\fifo0.fifo_store[27][0] ),
    .A1(_06033_),
    .S(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__clkbuf_1 _11463_ (.A(_06057_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _11464_ (.A0(\fifo0.fifo_store[27][1] ),
    .A1(_06037_),
    .S(_06056_),
    .X(_06058_));
 sky130_fd_sc_hd__clkbuf_1 _11465_ (.A(_06058_),
    .X(_01745_));
 sky130_fd_sc_hd__clkbuf_4 _11466_ (.A(_03875_),
    .X(_06059_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(\fifo0.fifo_store[27][2] ),
    .A1(_06059_),
    .S(_06056_),
    .X(_06060_));
 sky130_fd_sc_hd__clkbuf_1 _11468_ (.A(_06060_),
    .X(_01746_));
 sky130_fd_sc_hd__clkbuf_4 _11469_ (.A(_03878_),
    .X(_06061_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(\fifo0.fifo_store[27][3] ),
    .A1(_06061_),
    .S(_06056_),
    .X(_06062_));
 sky130_fd_sc_hd__clkbuf_1 _11471_ (.A(_06062_),
    .X(_01747_));
 sky130_fd_sc_hd__clkbuf_4 _11472_ (.A(_03881_),
    .X(_06063_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(\fifo0.fifo_store[27][4] ),
    .A1(_06063_),
    .S(_06056_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _11474_ (.A(_06064_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _11475_ (.A0(\fifo0.fifo_store[27][5] ),
    .A1(_05869_),
    .S(_06056_),
    .X(_06065_));
 sky130_fd_sc_hd__clkbuf_1 _11476_ (.A(_06065_),
    .X(_01749_));
 sky130_fd_sc_hd__clkbuf_4 _11477_ (.A(_03887_),
    .X(_06066_));
 sky130_fd_sc_hd__mux2_1 _11478_ (.A0(\fifo0.fifo_store[27][6] ),
    .A1(_06066_),
    .S(_06056_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_1 _11479_ (.A(_06067_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _11480_ (.A0(\fifo0.fifo_store[27][7] ),
    .A1(_05872_),
    .S(_06056_),
    .X(_06068_));
 sky130_fd_sc_hd__clkbuf_1 _11481_ (.A(_06068_),
    .X(_01751_));
 sky130_fd_sc_hd__clkbuf_4 _11482_ (.A(_03893_),
    .X(_06069_));
 sky130_fd_sc_hd__mux2_1 _11483_ (.A0(\fifo0.fifo_store[27][8] ),
    .A1(_06069_),
    .S(_06056_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_1 _11484_ (.A(_06070_),
    .X(_01752_));
 sky130_fd_sc_hd__clkbuf_4 _11485_ (.A(_03896_),
    .X(_06071_));
 sky130_fd_sc_hd__mux2_1 _11486_ (.A0(\fifo0.fifo_store[27][9] ),
    .A1(_06071_),
    .S(_06056_),
    .X(_06072_));
 sky130_fd_sc_hd__clkbuf_1 _11487_ (.A(_06072_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _11488_ (.A0(\fifo0.fifo_store[27][10] ),
    .A1(_05876_),
    .S(_06055_),
    .X(_06073_));
 sky130_fd_sc_hd__clkbuf_1 _11489_ (.A(_06073_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _11490_ (.A0(\fifo0.fifo_store[27][11] ),
    .A1(_05878_),
    .S(_06055_),
    .X(_06074_));
 sky130_fd_sc_hd__clkbuf_1 _11491_ (.A(_06074_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _11492_ (.A0(\fifo0.fifo_store[27][12] ),
    .A1(_06028_),
    .S(_06055_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _11493_ (.A(_06075_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(\fifo0.fifo_store[27][13] ),
    .A1(_06050_),
    .S(_06055_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_1 _11495_ (.A(_06076_),
    .X(_01757_));
 sky130_fd_sc_hd__clkbuf_4 _11496_ (.A(_03911_),
    .X(_06077_));
 sky130_fd_sc_hd__mux2_1 _11497_ (.A0(\fifo0.fifo_store[27][14] ),
    .A1(_06077_),
    .S(_06055_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _11498_ (.A(_06078_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _11499_ (.A0(\fifo0.fifo_store[27][15] ),
    .A1(_06053_),
    .S(_06055_),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_1 _11500_ (.A(_06079_),
    .X(_01759_));
 sky130_fd_sc_hd__nor2_8 _11501_ (.A(_03989_),
    .B(_05788_),
    .Y(_06080_));
 sky130_fd_sc_hd__buf_8 _11502_ (.A(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(\fifo0.fifo_store[26][0] ),
    .A1(_06033_),
    .S(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _11504_ (.A(_06082_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(\fifo0.fifo_store[26][1] ),
    .A1(_06037_),
    .S(_06081_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _11506_ (.A(_06083_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(\fifo0.fifo_store[26][2] ),
    .A1(_06059_),
    .S(_06081_),
    .X(_06084_));
 sky130_fd_sc_hd__clkbuf_1 _11508_ (.A(_06084_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(\fifo0.fifo_store[26][3] ),
    .A1(_06061_),
    .S(_06081_),
    .X(_06085_));
 sky130_fd_sc_hd__clkbuf_1 _11510_ (.A(_06085_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(\fifo0.fifo_store[26][4] ),
    .A1(_06063_),
    .S(_06081_),
    .X(_06086_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_06086_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(\fifo0.fifo_store[26][5] ),
    .A1(_05869_),
    .S(_06081_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _11514_ (.A(_06087_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\fifo0.fifo_store[26][6] ),
    .A1(_06066_),
    .S(_06081_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _11516_ (.A(_06088_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(\fifo0.fifo_store[26][7] ),
    .A1(_05872_),
    .S(_06081_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_1 _11518_ (.A(_06089_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(\fifo0.fifo_store[26][8] ),
    .A1(_06069_),
    .S(_06081_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _11520_ (.A(_06090_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(\fifo0.fifo_store[26][9] ),
    .A1(_06071_),
    .S(_06081_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _11522_ (.A(_06091_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(\fifo0.fifo_store[26][10] ),
    .A1(_05876_),
    .S(_06080_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _11524_ (.A(_06092_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _11525_ (.A0(\fifo0.fifo_store[26][11] ),
    .A1(_05878_),
    .S(_06080_),
    .X(_06093_));
 sky130_fd_sc_hd__clkbuf_1 _11526_ (.A(_06093_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(\fifo0.fifo_store[26][12] ),
    .A1(_06028_),
    .S(_06080_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _11528_ (.A(_06094_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _11529_ (.A0(\fifo0.fifo_store[26][13] ),
    .A1(_06050_),
    .S(_06080_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _11530_ (.A(_06095_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _11531_ (.A0(\fifo0.fifo_store[26][14] ),
    .A1(_06077_),
    .S(_06080_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _11532_ (.A(_06096_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _11533_ (.A0(\fifo0.fifo_store[26][15] ),
    .A1(_06053_),
    .S(_06080_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _11534_ (.A(_06097_),
    .X(_01775_));
 sky130_fd_sc_hd__nor2_8 _11535_ (.A(_04031_),
    .B(_05788_),
    .Y(_06098_));
 sky130_fd_sc_hd__buf_8 _11536_ (.A(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__mux2_1 _11537_ (.A0(\fifo0.fifo_store[25][0] ),
    .A1(\fifo0.fifo_data[0] ),
    .S(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _11538_ (.A(_06100_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _11539_ (.A0(\fifo0.fifo_store[25][1] ),
    .A1(\fifo0.fifo_data[1] ),
    .S(_06099_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _11540_ (.A(_06101_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _11541_ (.A0(\fifo0.fifo_store[25][2] ),
    .A1(\fifo0.fifo_data[2] ),
    .S(_06099_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _11542_ (.A(_06102_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _11543_ (.A0(\fifo0.fifo_store[25][3] ),
    .A1(\fifo0.fifo_data[3] ),
    .S(_06099_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_1 _11544_ (.A(_06103_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _11545_ (.A0(\fifo0.fifo_store[25][4] ),
    .A1(\fifo0.fifo_data[4] ),
    .S(_06099_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _11546_ (.A(_06104_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _11547_ (.A0(\fifo0.fifo_store[25][5] ),
    .A1(_05869_),
    .S(_06099_),
    .X(_06105_));
 sky130_fd_sc_hd__clkbuf_1 _11548_ (.A(_06105_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _11549_ (.A0(\fifo0.fifo_store[25][6] ),
    .A1(\fifo0.fifo_data[6] ),
    .S(_06099_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _11550_ (.A(_06106_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _11551_ (.A0(\fifo0.fifo_store[25][7] ),
    .A1(_05872_),
    .S(_06099_),
    .X(_06107_));
 sky130_fd_sc_hd__clkbuf_1 _11552_ (.A(_06107_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _11553_ (.A0(\fifo0.fifo_store[25][8] ),
    .A1(\fifo0.fifo_data[8] ),
    .S(_06099_),
    .X(_06108_));
 sky130_fd_sc_hd__clkbuf_1 _11554_ (.A(_06108_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _11555_ (.A0(\fifo0.fifo_store[25][9] ),
    .A1(\fifo0.fifo_data[9] ),
    .S(_06099_),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_1 _11556_ (.A(_06109_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _11557_ (.A0(\fifo0.fifo_store[25][10] ),
    .A1(_05876_),
    .S(_06098_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _11558_ (.A(_06110_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(\fifo0.fifo_store[25][11] ),
    .A1(_05878_),
    .S(_06098_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_1 _11560_ (.A(_06111_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(\fifo0.fifo_store[25][12] ),
    .A1(\fifo0.fifo_data[12] ),
    .S(_06098_),
    .X(_06112_));
 sky130_fd_sc_hd__clkbuf_1 _11562_ (.A(_06112_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(\fifo0.fifo_store[25][13] ),
    .A1(\fifo0.fifo_data[13] ),
    .S(_06098_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _11564_ (.A(_06113_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _11565_ (.A0(\fifo0.fifo_store[25][14] ),
    .A1(_06077_),
    .S(_06098_),
    .X(_06114_));
 sky130_fd_sc_hd__clkbuf_1 _11566_ (.A(_06114_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _11567_ (.A0(\fifo0.fifo_store[25][15] ),
    .A1(\fifo0.fifo_data[15] ),
    .S(_06098_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _11568_ (.A(_06115_),
    .X(_01791_));
 sky130_fd_sc_hd__nor2_8 _11569_ (.A(_03815_),
    .B(_05788_),
    .Y(_06116_));
 sky130_fd_sc_hd__buf_8 _11570_ (.A(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__mux2_1 _11571_ (.A0(\fifo0.fifo_store[24][0] ),
    .A1(_06033_),
    .S(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_1 _11572_ (.A(_06118_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\fifo0.fifo_store[24][1] ),
    .A1(_06037_),
    .S(_06117_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_1 _11574_ (.A(_06119_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(\fifo0.fifo_store[24][2] ),
    .A1(_06059_),
    .S(_06117_),
    .X(_06120_));
 sky130_fd_sc_hd__clkbuf_1 _11576_ (.A(_06120_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(\fifo0.fifo_store[24][3] ),
    .A1(_06061_),
    .S(_06117_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_1 _11578_ (.A(_06121_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _11579_ (.A0(\fifo0.fifo_store[24][4] ),
    .A1(_06063_),
    .S(_06117_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_1 _11580_ (.A(_06122_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_4 _11581_ (.A(_03838_),
    .X(_06123_));
 sky130_fd_sc_hd__mux2_1 _11582_ (.A0(\fifo0.fifo_store[24][5] ),
    .A1(_06123_),
    .S(_06117_),
    .X(_06124_));
 sky130_fd_sc_hd__clkbuf_1 _11583_ (.A(_06124_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _11584_ (.A0(\fifo0.fifo_store[24][6] ),
    .A1(_06066_),
    .S(_06117_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_1 _11585_ (.A(_06125_),
    .X(_01798_));
 sky130_fd_sc_hd__buf_4 _11586_ (.A(_03843_),
    .X(_06126_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(\fifo0.fifo_store[24][7] ),
    .A1(_06126_),
    .S(_06117_),
    .X(_06127_));
 sky130_fd_sc_hd__clkbuf_1 _11588_ (.A(_06127_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(\fifo0.fifo_store[24][8] ),
    .A1(_06069_),
    .S(_06117_),
    .X(_06128_));
 sky130_fd_sc_hd__clkbuf_1 _11590_ (.A(_06128_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(\fifo0.fifo_store[24][9] ),
    .A1(_06071_),
    .S(_06117_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_1 _11592_ (.A(_06129_),
    .X(_01801_));
 sky130_fd_sc_hd__buf_4 _11593_ (.A(_03850_),
    .X(_06130_));
 sky130_fd_sc_hd__mux2_1 _11594_ (.A0(\fifo0.fifo_store[24][10] ),
    .A1(_06130_),
    .S(_06116_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _11595_ (.A(_06131_),
    .X(_01802_));
 sky130_fd_sc_hd__buf_6 _11596_ (.A(_03853_),
    .X(_06132_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(\fifo0.fifo_store[24][11] ),
    .A1(_06132_),
    .S(_06116_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_1 _11598_ (.A(_06133_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _11599_ (.A0(\fifo0.fifo_store[24][12] ),
    .A1(_06028_),
    .S(_06116_),
    .X(_06134_));
 sky130_fd_sc_hd__clkbuf_1 _11600_ (.A(_06134_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _11601_ (.A0(\fifo0.fifo_store[24][13] ),
    .A1(_06050_),
    .S(_06116_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_1 _11602_ (.A(_06135_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _11603_ (.A0(\fifo0.fifo_store[24][14] ),
    .A1(_06077_),
    .S(_06116_),
    .X(_06136_));
 sky130_fd_sc_hd__clkbuf_1 _11604_ (.A(_06136_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(\fifo0.fifo_store[24][15] ),
    .A1(_06053_),
    .S(_06116_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_1 _11606_ (.A(_06137_),
    .X(_01807_));
 sky130_fd_sc_hd__nor2_8 _11607_ (.A(_03919_),
    .B(_05995_),
    .Y(_06138_));
 sky130_fd_sc_hd__buf_8 _11608_ (.A(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__mux2_1 _11609_ (.A0(\fifo0.fifo_store[23][0] ),
    .A1(_06033_),
    .S(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__clkbuf_1 _11610_ (.A(_06140_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(\fifo0.fifo_store[23][1] ),
    .A1(_06037_),
    .S(_06139_),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_1 _11612_ (.A(_06141_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(\fifo0.fifo_store[23][2] ),
    .A1(_06059_),
    .S(_06139_),
    .X(_06142_));
 sky130_fd_sc_hd__clkbuf_1 _11614_ (.A(_06142_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(\fifo0.fifo_store[23][3] ),
    .A1(_06061_),
    .S(_06139_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _11616_ (.A(_06143_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\fifo0.fifo_store[23][4] ),
    .A1(_06063_),
    .S(_06139_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _11618_ (.A(_06144_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(\fifo0.fifo_store[23][5] ),
    .A1(_06123_),
    .S(_06139_),
    .X(_06145_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_06145_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _11621_ (.A0(\fifo0.fifo_store[23][6] ),
    .A1(_06066_),
    .S(_06139_),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_1 _11622_ (.A(_06146_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(\fifo0.fifo_store[23][7] ),
    .A1(_06126_),
    .S(_06139_),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _11624_ (.A(_06147_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _11625_ (.A0(\fifo0.fifo_store[23][8] ),
    .A1(_06069_),
    .S(_06139_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _11626_ (.A(_06148_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(\fifo0.fifo_store[23][9] ),
    .A1(_06071_),
    .S(_06139_),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _11628_ (.A(_06149_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _11629_ (.A0(\fifo0.fifo_store[23][10] ),
    .A1(_06130_),
    .S(_06138_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _11630_ (.A(_06150_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(\fifo0.fifo_store[23][11] ),
    .A1(_06132_),
    .S(_06138_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _11632_ (.A(_06151_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _11633_ (.A0(\fifo0.fifo_store[23][12] ),
    .A1(_06028_),
    .S(_06138_),
    .X(_06152_));
 sky130_fd_sc_hd__clkbuf_1 _11634_ (.A(_06152_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _11635_ (.A0(\fifo0.fifo_store[23][13] ),
    .A1(_06050_),
    .S(_06138_),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_1 _11636_ (.A(_06153_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(\fifo0.fifo_store[23][14] ),
    .A1(_06077_),
    .S(_06138_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_06154_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(\fifo0.fifo_store[23][15] ),
    .A1(_06053_),
    .S(_06138_),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _11640_ (.A(_06155_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _11641_ (.A(_03943_),
    .B(_05995_),
    .X(_06156_));
 sky130_fd_sc_hd__buf_4 _11642_ (.A(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__buf_8 _11643_ (.A(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__mux2_1 _11644_ (.A0(_04885_),
    .A1(\fifo0.fifo_store[22][0] ),
    .S(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _11645_ (.A(_06159_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(_04890_),
    .A1(\fifo0.fifo_store[22][1] ),
    .S(_06158_),
    .X(_06160_));
 sky130_fd_sc_hd__clkbuf_1 _11647_ (.A(_06160_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(_04892_),
    .A1(\fifo0.fifo_store[22][2] ),
    .S(_06158_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _11649_ (.A(_06161_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _11650_ (.A0(_04894_),
    .A1(\fifo0.fifo_store[22][3] ),
    .S(_06158_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _11651_ (.A(_06162_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _11652_ (.A0(_04896_),
    .A1(\fifo0.fifo_store[22][4] ),
    .S(_06158_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _11653_ (.A(_06163_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(_04898_),
    .A1(\fifo0.fifo_store[22][5] ),
    .S(_06158_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _11655_ (.A(_06164_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(_04900_),
    .A1(\fifo0.fifo_store[22][6] ),
    .S(_06158_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _11657_ (.A(_06165_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(_04902_),
    .A1(\fifo0.fifo_store[22][7] ),
    .S(_06158_),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _11659_ (.A(_06166_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(_04904_),
    .A1(\fifo0.fifo_store[22][8] ),
    .S(_06158_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _11661_ (.A(_06167_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(_04906_),
    .A1(\fifo0.fifo_store[22][9] ),
    .S(_06158_),
    .X(_06168_));
 sky130_fd_sc_hd__clkbuf_1 _11663_ (.A(_06168_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(_04908_),
    .A1(\fifo0.fifo_store[22][10] ),
    .S(_06157_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _11665_ (.A(_06169_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(_04910_),
    .A1(\fifo0.fifo_store[22][11] ),
    .S(_06157_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _11667_ (.A(_06170_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(_04912_),
    .A1(\fifo0.fifo_store[22][12] ),
    .S(_06157_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _11669_ (.A(_06171_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(_04914_),
    .A1(\fifo0.fifo_store[22][13] ),
    .S(_06157_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _11671_ (.A(_06172_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(_04916_),
    .A1(\fifo0.fifo_store[22][14] ),
    .S(_06157_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _11673_ (.A(_06173_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(_04918_),
    .A1(\fifo0.fifo_store[22][15] ),
    .S(_06157_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _11675_ (.A(_06174_),
    .X(_01839_));
 sky130_fd_sc_hd__nor2_8 _11676_ (.A(_03964_),
    .B(_05995_),
    .Y(_06175_));
 sky130_fd_sc_hd__clkbuf_16 _11677_ (.A(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(\fifo0.fifo_store[21][0] ),
    .A1(_06033_),
    .S(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _11679_ (.A(_06177_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(\fifo0.fifo_store[21][1] ),
    .A1(_06037_),
    .S(_06176_),
    .X(_06178_));
 sky130_fd_sc_hd__clkbuf_1 _11681_ (.A(_06178_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _11682_ (.A0(\fifo0.fifo_store[21][2] ),
    .A1(_06059_),
    .S(_06176_),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_1 _11683_ (.A(_06179_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(\fifo0.fifo_store[21][3] ),
    .A1(_06061_),
    .S(_06176_),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_1 _11685_ (.A(_06180_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(\fifo0.fifo_store[21][4] ),
    .A1(_06063_),
    .S(_06176_),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _11687_ (.A(_06181_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(\fifo0.fifo_store[21][5] ),
    .A1(_06123_),
    .S(_06176_),
    .X(_06182_));
 sky130_fd_sc_hd__clkbuf_1 _11689_ (.A(_06182_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(\fifo0.fifo_store[21][6] ),
    .A1(_06066_),
    .S(_06176_),
    .X(_06183_));
 sky130_fd_sc_hd__clkbuf_1 _11691_ (.A(_06183_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(\fifo0.fifo_store[21][7] ),
    .A1(_06126_),
    .S(_06176_),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_06184_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(\fifo0.fifo_store[21][8] ),
    .A1(_06069_),
    .S(_06176_),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_06185_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(\fifo0.fifo_store[21][9] ),
    .A1(_06071_),
    .S(_06176_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_06186_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(\fifo0.fifo_store[21][10] ),
    .A1(_06130_),
    .S(_06175_),
    .X(_06187_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_06187_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\fifo0.fifo_store[21][11] ),
    .A1(_06132_),
    .S(_06175_),
    .X(_06188_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_06188_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\fifo0.fifo_store[21][12] ),
    .A1(_06028_),
    .S(_06175_),
    .X(_06189_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_06189_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(\fifo0.fifo_store[21][13] ),
    .A1(_06050_),
    .S(_06175_),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_1 _11705_ (.A(_06190_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(\fifo0.fifo_store[21][14] ),
    .A1(_06077_),
    .S(_06175_),
    .X(_06191_));
 sky130_fd_sc_hd__clkbuf_1 _11707_ (.A(_06191_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(\fifo0.fifo_store[21][15] ),
    .A1(_06053_),
    .S(_06175_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _11709_ (.A(_06192_),
    .X(_01855_));
 sky130_fd_sc_hd__nor2_8 _11710_ (.A(_04010_),
    .B(_05995_),
    .Y(_06193_));
 sky130_fd_sc_hd__clkbuf_16 _11711_ (.A(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(\fifo0.fifo_store[20][0] ),
    .A1(_06033_),
    .S(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _11713_ (.A(_06195_),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(\fifo0.fifo_store[20][1] ),
    .A1(_06037_),
    .S(_06194_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_1 _11715_ (.A(_06196_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _11716_ (.A0(\fifo0.fifo_store[20][2] ),
    .A1(_06059_),
    .S(_06194_),
    .X(_06197_));
 sky130_fd_sc_hd__clkbuf_1 _11717_ (.A(_06197_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(\fifo0.fifo_store[20][3] ),
    .A1(_06061_),
    .S(_06194_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _11719_ (.A(_06198_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(\fifo0.fifo_store[20][4] ),
    .A1(_06063_),
    .S(_06194_),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_1 _11721_ (.A(_06199_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _11722_ (.A0(\fifo0.fifo_store[20][5] ),
    .A1(_06123_),
    .S(_06194_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_1 _11723_ (.A(_06200_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(\fifo0.fifo_store[20][6] ),
    .A1(_06066_),
    .S(_06194_),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_1 _11725_ (.A(_06201_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(\fifo0.fifo_store[20][7] ),
    .A1(_06126_),
    .S(_06194_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _11727_ (.A(_06202_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(\fifo0.fifo_store[20][8] ),
    .A1(_06069_),
    .S(_06194_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_1 _11729_ (.A(_06203_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(\fifo0.fifo_store[20][9] ),
    .A1(_06071_),
    .S(_06194_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_06204_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(\fifo0.fifo_store[20][10] ),
    .A1(_06130_),
    .S(_06193_),
    .X(_06205_));
 sky130_fd_sc_hd__clkbuf_1 _11733_ (.A(_06205_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\fifo0.fifo_store[20][11] ),
    .A1(_06132_),
    .S(_06193_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_1 _11735_ (.A(_06206_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\fifo0.fifo_store[20][12] ),
    .A1(_06028_),
    .S(_06193_),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_06207_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(\fifo0.fifo_store[20][13] ),
    .A1(_06050_),
    .S(_06193_),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_1 _11739_ (.A(_06208_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(\fifo0.fifo_store[20][14] ),
    .A1(_06077_),
    .S(_06193_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _11741_ (.A(_06209_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\fifo0.fifo_store[20][15] ),
    .A1(_06053_),
    .S(_06193_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _11743_ (.A(_06210_),
    .X(_01871_));
 sky130_fd_sc_hd__nor2_8 _11744_ (.A(_03814_),
    .B(_04032_),
    .Y(_06211_));
 sky130_fd_sc_hd__buf_6 _11745_ (.A(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(\fifo0.fifo_store[1][0] ),
    .A1(_06033_),
    .S(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _11747_ (.A(_06213_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(\fifo0.fifo_store[1][1] ),
    .A1(_06037_),
    .S(_06212_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_06214_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(\fifo0.fifo_store[1][2] ),
    .A1(_06059_),
    .S(_06212_),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_1 _11751_ (.A(_06215_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(\fifo0.fifo_store[1][3] ),
    .A1(_06061_),
    .S(_06212_),
    .X(_06216_));
 sky130_fd_sc_hd__clkbuf_1 _11753_ (.A(_06216_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(\fifo0.fifo_store[1][4] ),
    .A1(_06063_),
    .S(_06212_),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _11755_ (.A(_06217_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(\fifo0.fifo_store[1][5] ),
    .A1(_06123_),
    .S(_06212_),
    .X(_06218_));
 sky130_fd_sc_hd__clkbuf_1 _11757_ (.A(_06218_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(\fifo0.fifo_store[1][6] ),
    .A1(_06066_),
    .S(_06212_),
    .X(_06219_));
 sky130_fd_sc_hd__clkbuf_1 _11759_ (.A(_06219_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(\fifo0.fifo_store[1][7] ),
    .A1(_06126_),
    .S(_06212_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _11761_ (.A(_06220_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(\fifo0.fifo_store[1][8] ),
    .A1(_06069_),
    .S(_06212_),
    .X(_06221_));
 sky130_fd_sc_hd__clkbuf_1 _11763_ (.A(_06221_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(\fifo0.fifo_store[1][9] ),
    .A1(_06071_),
    .S(_06212_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _11765_ (.A(_06222_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(\fifo0.fifo_store[1][10] ),
    .A1(_06130_),
    .S(_06211_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _11767_ (.A(_06223_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(\fifo0.fifo_store[1][11] ),
    .A1(_06132_),
    .S(_06211_),
    .X(_06224_));
 sky130_fd_sc_hd__clkbuf_1 _11769_ (.A(_06224_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(\fifo0.fifo_store[1][12] ),
    .A1(_06028_),
    .S(_06211_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _11771_ (.A(_06225_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(\fifo0.fifo_store[1][13] ),
    .A1(_06050_),
    .S(_06211_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _11773_ (.A(_06226_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(\fifo0.fifo_store[1][14] ),
    .A1(_06077_),
    .S(_06211_),
    .X(_06227_));
 sky130_fd_sc_hd__clkbuf_1 _11775_ (.A(_06227_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(\fifo0.fifo_store[1][15] ),
    .A1(_06053_),
    .S(_06211_),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_1 _11777_ (.A(_06228_),
    .X(_01887_));
 sky130_fd_sc_hd__and2_1 _11778_ (.A(_05916_),
    .B(\fifo0.fifo_data_del1[0] ),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _11779_ (.A(_06229_),
    .X(_01888_));
 sky130_fd_sc_hd__and2_1 _11780_ (.A(_05916_),
    .B(\fifo0.fifo_data_del1[1] ),
    .X(_06230_));
 sky130_fd_sc_hd__clkbuf_1 _11781_ (.A(_06230_),
    .X(_01889_));
 sky130_fd_sc_hd__and2_1 _11782_ (.A(_05916_),
    .B(\fifo0.fifo_data_del1[2] ),
    .X(_06231_));
 sky130_fd_sc_hd__clkbuf_1 _11783_ (.A(_06231_),
    .X(_01890_));
 sky130_fd_sc_hd__clkbuf_4 _11784_ (.A(net21),
    .X(_06232_));
 sky130_fd_sc_hd__and2_1 _11785_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[3] ),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _11786_ (.A(_06233_),
    .X(_01891_));
 sky130_fd_sc_hd__and2_1 _11787_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[4] ),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_1 _11788_ (.A(_06234_),
    .X(_01892_));
 sky130_fd_sc_hd__and2_1 _11789_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[5] ),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_1 _11790_ (.A(_06235_),
    .X(_01893_));
 sky130_fd_sc_hd__and2_1 _11791_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[6] ),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _11792_ (.A(_06236_),
    .X(_01894_));
 sky130_fd_sc_hd__and2_1 _11793_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[7] ),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _11794_ (.A(_06237_),
    .X(_01895_));
 sky130_fd_sc_hd__and2_1 _11795_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[8] ),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _11796_ (.A(_06238_),
    .X(_01896_));
 sky130_fd_sc_hd__and2_1 _11797_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[9] ),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _11798_ (.A(_06239_),
    .X(_01897_));
 sky130_fd_sc_hd__and2_1 _11799_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[10] ),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_1 _11800_ (.A(_06240_),
    .X(_01898_));
 sky130_fd_sc_hd__and2_1 _11801_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[11] ),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _11802_ (.A(_06241_),
    .X(_01899_));
 sky130_fd_sc_hd__and2_1 _11803_ (.A(_06232_),
    .B(\fifo0.fifo_data_del1[12] ),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_1 _11804_ (.A(_06242_),
    .X(_01900_));
 sky130_fd_sc_hd__and2_1 _11805_ (.A(_05902_),
    .B(\fifo0.fifo_data_del1[13] ),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _11806_ (.A(_06243_),
    .X(_01901_));
 sky130_fd_sc_hd__and2_1 _11807_ (.A(_05902_),
    .B(\fifo0.fifo_data_del1[14] ),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _11808_ (.A(_06244_),
    .X(_01902_));
 sky130_fd_sc_hd__and2_1 _11809_ (.A(_05902_),
    .B(\fifo0.fifo_data_del1[15] ),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _11810_ (.A(_06245_),
    .X(_01903_));
 sky130_fd_sc_hd__nor2_8 _11811_ (.A(_03919_),
    .B(_03941_),
    .Y(_06246_));
 sky130_fd_sc_hd__buf_6 _11812_ (.A(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(\fifo0.fifo_store[79][0] ),
    .A1(_06033_),
    .S(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _11814_ (.A(_06248_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(\fifo0.fifo_store[79][1] ),
    .A1(_06037_),
    .S(_06247_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _11816_ (.A(_06249_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(\fifo0.fifo_store[79][2] ),
    .A1(_06059_),
    .S(_06247_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _11818_ (.A(_06250_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(\fifo0.fifo_store[79][3] ),
    .A1(_06061_),
    .S(_06247_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _11820_ (.A(_06251_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(\fifo0.fifo_store[79][4] ),
    .A1(_06063_),
    .S(_06247_),
    .X(_06252_));
 sky130_fd_sc_hd__clkbuf_1 _11822_ (.A(_06252_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(\fifo0.fifo_store[79][5] ),
    .A1(_06123_),
    .S(_06247_),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_1 _11824_ (.A(_06253_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(\fifo0.fifo_store[79][6] ),
    .A1(_06066_),
    .S(_06247_),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_1 _11826_ (.A(_06254_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(\fifo0.fifo_store[79][7] ),
    .A1(_06126_),
    .S(_06247_),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_1 _11828_ (.A(_06255_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _11829_ (.A0(\fifo0.fifo_store[79][8] ),
    .A1(_06069_),
    .S(_06247_),
    .X(_06256_));
 sky130_fd_sc_hd__clkbuf_1 _11830_ (.A(_06256_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(\fifo0.fifo_store[79][9] ),
    .A1(_06071_),
    .S(_06247_),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_1 _11832_ (.A(_06257_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(\fifo0.fifo_store[79][10] ),
    .A1(_06130_),
    .S(_06246_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _11834_ (.A(_06258_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(\fifo0.fifo_store[79][11] ),
    .A1(_06132_),
    .S(_06246_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _11836_ (.A(_06259_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(\fifo0.fifo_store[79][12] ),
    .A1(_06028_),
    .S(_06246_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _11838_ (.A(_06260_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _11839_ (.A0(\fifo0.fifo_store[79][13] ),
    .A1(_06050_),
    .S(_06246_),
    .X(_06261_));
 sky130_fd_sc_hd__clkbuf_1 _11840_ (.A(_06261_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _11841_ (.A0(\fifo0.fifo_store[79][14] ),
    .A1(_06077_),
    .S(_06246_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _11842_ (.A(_06262_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(\fifo0.fifo_store[79][15] ),
    .A1(_06053_),
    .S(_06246_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _11844_ (.A(_06263_),
    .X(_01919_));
 sky130_fd_sc_hd__nor2_8 _11845_ (.A(_03989_),
    .B(_05995_),
    .Y(_06264_));
 sky130_fd_sc_hd__buf_8 _11846_ (.A(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\fifo0.fifo_store[18][0] ),
    .A1(_06033_),
    .S(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _11848_ (.A(_06266_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(\fifo0.fifo_store[18][1] ),
    .A1(_06037_),
    .S(_06265_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _11850_ (.A(_06267_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(\fifo0.fifo_store[18][2] ),
    .A1(_06059_),
    .S(_06265_),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _11852_ (.A(_06268_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(\fifo0.fifo_store[18][3] ),
    .A1(_06061_),
    .S(_06265_),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_1 _11854_ (.A(_06269_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(\fifo0.fifo_store[18][4] ),
    .A1(_06063_),
    .S(_06265_),
    .X(_06270_));
 sky130_fd_sc_hd__clkbuf_1 _11856_ (.A(_06270_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(\fifo0.fifo_store[18][5] ),
    .A1(_06123_),
    .S(_06265_),
    .X(_06271_));
 sky130_fd_sc_hd__clkbuf_1 _11858_ (.A(_06271_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\fifo0.fifo_store[18][6] ),
    .A1(_06066_),
    .S(_06265_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _11860_ (.A(_06272_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\fifo0.fifo_store[18][7] ),
    .A1(_06126_),
    .S(_06265_),
    .X(_06273_));
 sky130_fd_sc_hd__clkbuf_1 _11862_ (.A(_06273_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(\fifo0.fifo_store[18][8] ),
    .A1(_06069_),
    .S(_06265_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_06274_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\fifo0.fifo_store[18][9] ),
    .A1(_06071_),
    .S(_06265_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_06275_),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\fifo0.fifo_store[18][10] ),
    .A1(_06130_),
    .S(_06264_),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_06276_),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\fifo0.fifo_store[18][11] ),
    .A1(_06132_),
    .S(_06264_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_06277_),
    .X(_01931_));
 sky130_fd_sc_hd__buf_6 _11871_ (.A(_03855_),
    .X(_06278_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(\fifo0.fifo_store[18][12] ),
    .A1(_06278_),
    .S(_06264_),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _11873_ (.A(_06279_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(\fifo0.fifo_store[18][13] ),
    .A1(_06050_),
    .S(_06264_),
    .X(_06280_));
 sky130_fd_sc_hd__clkbuf_1 _11875_ (.A(_06280_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\fifo0.fifo_store[18][14] ),
    .A1(_06077_),
    .S(_06264_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _11877_ (.A(_06281_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(\fifo0.fifo_store[18][15] ),
    .A1(_06053_),
    .S(_06264_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(_06282_),
    .X(_01935_));
 sky130_fd_sc_hd__buf_4 _11880_ (.A(_03820_),
    .X(_06283_));
 sky130_fd_sc_hd__nor2_8 _11881_ (.A(_04010_),
    .B(_04356_),
    .Y(_06284_));
 sky130_fd_sc_hd__buf_8 _11882_ (.A(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_1 _11883_ (.A0(\fifo0.fifo_store[12][0] ),
    .A1(_06283_),
    .S(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _11884_ (.A(_06286_),
    .X(_01936_));
 sky130_fd_sc_hd__buf_4 _11885_ (.A(_03828_),
    .X(_06287_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\fifo0.fifo_store[12][1] ),
    .A1(_06287_),
    .S(_06285_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _11887_ (.A(_06288_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\fifo0.fifo_store[12][2] ),
    .A1(_06059_),
    .S(_06285_),
    .X(_06289_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_06289_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(\fifo0.fifo_store[12][3] ),
    .A1(_06061_),
    .S(_06285_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _11891_ (.A(_06290_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(\fifo0.fifo_store[12][4] ),
    .A1(_06063_),
    .S(_06285_),
    .X(_06291_));
 sky130_fd_sc_hd__clkbuf_1 _11893_ (.A(_06291_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(\fifo0.fifo_store[12][5] ),
    .A1(_06123_),
    .S(_06285_),
    .X(_06292_));
 sky130_fd_sc_hd__clkbuf_1 _11895_ (.A(_06292_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(\fifo0.fifo_store[12][6] ),
    .A1(_06066_),
    .S(_06285_),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _11897_ (.A(_06293_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(\fifo0.fifo_store[12][7] ),
    .A1(_06126_),
    .S(_06285_),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _11899_ (.A(_06294_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(\fifo0.fifo_store[12][8] ),
    .A1(_06069_),
    .S(_06285_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_1 _11901_ (.A(_06295_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(\fifo0.fifo_store[12][9] ),
    .A1(_06071_),
    .S(_06285_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _11903_ (.A(_06296_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(\fifo0.fifo_store[12][10] ),
    .A1(_06130_),
    .S(_06284_),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_1 _11905_ (.A(_06297_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(\fifo0.fifo_store[12][11] ),
    .A1(_06132_),
    .S(_06284_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_1 _11907_ (.A(_06298_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(\fifo0.fifo_store[12][12] ),
    .A1(_06278_),
    .S(_06284_),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _11909_ (.A(_06299_),
    .X(_01948_));
 sky130_fd_sc_hd__buf_6 _11910_ (.A(_03857_),
    .X(_06300_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(\fifo0.fifo_store[12][13] ),
    .A1(_06300_),
    .S(_06284_),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _11912_ (.A(_06301_),
    .X(_01949_));
 sky130_fd_sc_hd__buf_8 _11913_ (.A(_03859_),
    .X(_06302_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(\fifo0.fifo_store[12][14] ),
    .A1(_06302_),
    .S(_06284_),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _11915_ (.A(_06303_),
    .X(_01950_));
 sky130_fd_sc_hd__buf_6 _11916_ (.A(_03861_),
    .X(_06304_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\fifo0.fifo_store[12][15] ),
    .A1(_06304_),
    .S(_06284_),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _11918_ (.A(_06305_),
    .X(_01951_));
 sky130_fd_sc_hd__nor2_8 _11919_ (.A(_04052_),
    .B(_05995_),
    .Y(_06306_));
 sky130_fd_sc_hd__buf_8 _11920_ (.A(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(\fifo0.fifo_store[19][0] ),
    .A1(_06283_),
    .S(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(_06308_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(\fifo0.fifo_store[19][1] ),
    .A1(_06287_),
    .S(_06307_),
    .X(_06309_));
 sky130_fd_sc_hd__clkbuf_1 _11924_ (.A(_06309_),
    .X(_01953_));
 sky130_fd_sc_hd__buf_6 _11925_ (.A(_03875_),
    .X(_06310_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(\fifo0.fifo_store[19][2] ),
    .A1(_06310_),
    .S(_06307_),
    .X(_06311_));
 sky130_fd_sc_hd__clkbuf_1 _11927_ (.A(_06311_),
    .X(_01954_));
 sky130_fd_sc_hd__buf_4 _11928_ (.A(_03878_),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(\fifo0.fifo_store[19][3] ),
    .A1(_06312_),
    .S(_06307_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_1 _11930_ (.A(_06313_),
    .X(_01955_));
 sky130_fd_sc_hd__clkbuf_8 _11931_ (.A(_03881_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _11932_ (.A0(\fifo0.fifo_store[19][4] ),
    .A1(_06314_),
    .S(_06307_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _11933_ (.A(_06315_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(\fifo0.fifo_store[19][5] ),
    .A1(_06123_),
    .S(_06307_),
    .X(_06316_));
 sky130_fd_sc_hd__clkbuf_1 _11935_ (.A(_06316_),
    .X(_01957_));
 sky130_fd_sc_hd__buf_6 _11936_ (.A(_03887_),
    .X(_06317_));
 sky130_fd_sc_hd__mux2_1 _11937_ (.A0(\fifo0.fifo_store[19][6] ),
    .A1(_06317_),
    .S(_06307_),
    .X(_06318_));
 sky130_fd_sc_hd__clkbuf_1 _11938_ (.A(_06318_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _11939_ (.A0(\fifo0.fifo_store[19][7] ),
    .A1(_06126_),
    .S(_06307_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _11940_ (.A(_06319_),
    .X(_01959_));
 sky130_fd_sc_hd__buf_6 _11941_ (.A(_03893_),
    .X(_06320_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\fifo0.fifo_store[19][8] ),
    .A1(_06320_),
    .S(_06307_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _11943_ (.A(_06321_),
    .X(_01960_));
 sky130_fd_sc_hd__buf_4 _11944_ (.A(_03896_),
    .X(_06322_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(\fifo0.fifo_store[19][9] ),
    .A1(_06322_),
    .S(_06307_),
    .X(_06323_));
 sky130_fd_sc_hd__clkbuf_1 _11946_ (.A(_06323_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(\fifo0.fifo_store[19][10] ),
    .A1(_06130_),
    .S(_06306_),
    .X(_06324_));
 sky130_fd_sc_hd__clkbuf_1 _11948_ (.A(_06324_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(\fifo0.fifo_store[19][11] ),
    .A1(_06132_),
    .S(_06306_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _11950_ (.A(_06325_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(\fifo0.fifo_store[19][12] ),
    .A1(_06278_),
    .S(_06306_),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_1 _11952_ (.A(_06326_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(\fifo0.fifo_store[19][13] ),
    .A1(_06300_),
    .S(_06306_),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _11954_ (.A(_06327_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(\fifo0.fifo_store[19][14] ),
    .A1(_06302_),
    .S(_06306_),
    .X(_06328_));
 sky130_fd_sc_hd__clkbuf_1 _11956_ (.A(_06328_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(\fifo0.fifo_store[19][15] ),
    .A1(_06304_),
    .S(_06306_),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _11958_ (.A(_06329_),
    .X(_01967_));
 sky130_fd_sc_hd__nor2_8 _11959_ (.A(_03919_),
    .B(_04376_),
    .Y(_06330_));
 sky130_fd_sc_hd__buf_6 _11960_ (.A(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(\fifo0.fifo_store[127][0] ),
    .A1(_06283_),
    .S(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_06332_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(\fifo0.fifo_store[127][1] ),
    .A1(_06287_),
    .S(_06331_),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_06333_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(\fifo0.fifo_store[127][2] ),
    .A1(_06310_),
    .S(_06331_),
    .X(_06334_));
 sky130_fd_sc_hd__clkbuf_1 _11966_ (.A(_06334_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(\fifo0.fifo_store[127][3] ),
    .A1(_06312_),
    .S(_06331_),
    .X(_06335_));
 sky130_fd_sc_hd__clkbuf_1 _11968_ (.A(_06335_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(\fifo0.fifo_store[127][4] ),
    .A1(_06314_),
    .S(_06331_),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _11970_ (.A(_06336_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(\fifo0.fifo_store[127][5] ),
    .A1(_06123_),
    .S(_06331_),
    .X(_06337_));
 sky130_fd_sc_hd__clkbuf_1 _11972_ (.A(_06337_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(\fifo0.fifo_store[127][6] ),
    .A1(_06317_),
    .S(_06331_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_1 _11974_ (.A(_06338_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _11975_ (.A0(\fifo0.fifo_store[127][7] ),
    .A1(_06126_),
    .S(_06331_),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _11976_ (.A(_06339_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(\fifo0.fifo_store[127][8] ),
    .A1(_06320_),
    .S(_06331_),
    .X(_06340_));
 sky130_fd_sc_hd__clkbuf_1 _11978_ (.A(_06340_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(\fifo0.fifo_store[127][9] ),
    .A1(_06322_),
    .S(_06331_),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_1 _11980_ (.A(_06341_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(\fifo0.fifo_store[127][10] ),
    .A1(_06130_),
    .S(_06330_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_1 _11982_ (.A(_06342_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(\fifo0.fifo_store[127][11] ),
    .A1(_06132_),
    .S(_06330_),
    .X(_06343_));
 sky130_fd_sc_hd__clkbuf_1 _11984_ (.A(_06343_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(\fifo0.fifo_store[127][12] ),
    .A1(_06278_),
    .S(_06330_),
    .X(_06344_));
 sky130_fd_sc_hd__clkbuf_1 _11986_ (.A(_06344_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(\fifo0.fifo_store[127][13] ),
    .A1(_06300_),
    .S(_06330_),
    .X(_06345_));
 sky130_fd_sc_hd__clkbuf_1 _11988_ (.A(_06345_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\fifo0.fifo_store[127][14] ),
    .A1(_06302_),
    .S(_06330_),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_06346_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\fifo0.fifo_store[127][15] ),
    .A1(_06304_),
    .S(_06330_),
    .X(_06347_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_06347_),
    .X(_01983_));
 sky130_fd_sc_hd__clkbuf_4 _11993_ (.A(net18),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_4 _11994_ (.A(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a21oi_1 _11995_ (.A1(_06349_),
    .A2(\dsmod0.mod2_ctr[0] ),
    .B1(_05924_),
    .Y(_06350_));
 sky130_fd_sc_hd__o21a_1 _11996_ (.A1(_06349_),
    .A2(\dsmod0.mod2_ctr[0] ),
    .B1(_06350_),
    .X(_01984_));
 sky130_fd_sc_hd__a21oi_1 _11997_ (.A1(_06349_),
    .A2(\dsmod0.mod2_ctr[0] ),
    .B1(\dsmod0.mod2_ctr[1] ),
    .Y(_06351_));
 sky130_fd_sc_hd__a31o_1 _11998_ (.A1(_06349_),
    .A2(\dsmod0.mod2_ctr[1] ),
    .A3(\dsmod0.mod2_ctr[0] ),
    .B1(_05924_),
    .X(_06352_));
 sky130_fd_sc_hd__nor2_1 _11999_ (.A(_06351_),
    .B(_06352_),
    .Y(_01985_));
 sky130_fd_sc_hd__clkbuf_4 _12000_ (.A(net30),
    .X(_06353_));
 sky130_fd_sc_hd__clkbuf_4 _12001_ (.A(net33),
    .X(_06354_));
 sky130_fd_sc_hd__and4_1 _12002_ (.A(net31),
    .B(_06353_),
    .C(_06354_),
    .D(net32),
    .X(_06355_));
 sky130_fd_sc_hd__buf_2 _12003_ (.A(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__clkinv_4 _12004_ (.A(net23),
    .Y(_06357_));
 sky130_fd_sc_hd__clkbuf_4 _12005_ (.A(\sinegen0.read_ptr[4] ),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_4 _12006_ (.A(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__xnor2_2 _12007_ (.A(\sinegen0.read_ptr[1] ),
    .B(\sinegen0.read_ptr[0] ),
    .Y(_06360_));
 sky130_fd_sc_hd__clkbuf_4 _12008_ (.A(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__buf_2 _12009_ (.A(\sinegen0.read_ptr[3] ),
    .X(_06362_));
 sky130_fd_sc_hd__clkbuf_4 _12010_ (.A(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_4 _12011_ (.A(\sinegen0.read_ptr[1] ),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_4 _12012_ (.A(\sinegen0.read_ptr[0] ),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_4 _12013_ (.A(\sinegen0.read_ptr[2] ),
    .X(_06366_));
 sky130_fd_sc_hd__o21a_2 _12014_ (.A1(_06364_),
    .A2(_06365_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor2_1 _12015_ (.A(_06363_),
    .B(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__clkinv_2 _12016_ (.A(\sinegen0.read_ptr[5] ),
    .Y(_06369_));
 sky130_fd_sc_hd__clkbuf_4 _12017_ (.A(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__o211a_1 _12018_ (.A1(_06359_),
    .A2(_06361_),
    .B1(_06368_),
    .C1(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__nand3_1 _12019_ (.A(_06362_),
    .B(_06366_),
    .C(_06364_),
    .Y(_06372_));
 sky130_fd_sc_hd__buf_2 _12020_ (.A(\sinegen0.read_ptr[4] ),
    .X(_06373_));
 sky130_fd_sc_hd__or2_2 _12021_ (.A(\sinegen0.read_ptr[5] ),
    .B(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__nor2_1 _12022_ (.A(_06372_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__buf_4 _12023_ (.A(\sinegen0.read_ptr[3] ),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_4 _12024_ (.A(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_4 _12025_ (.A(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_4 _12026_ (.A(\sinegen0.read_ptr[1] ),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_4 _12027_ (.A(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__and2_1 _12028_ (.A(\sinegen0.read_ptr[2] ),
    .B(\sinegen0.read_ptr[0] ),
    .X(_06381_));
 sky130_fd_sc_hd__buf_2 _12029_ (.A(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__nand2_1 _12030_ (.A(_06380_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__or3b_4 _12031_ (.A(\sinegen0.read_ptr[2] ),
    .B(\sinegen0.read_ptr[0] ),
    .C_N(\sinegen0.read_ptr[1] ),
    .X(_06384_));
 sky130_fd_sc_hd__or2_1 _12032_ (.A(\sinegen0.read_ptr[2] ),
    .B(\sinegen0.read_ptr[1] ),
    .X(_06385_));
 sky130_fd_sc_hd__buf_2 _12033_ (.A(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__nor2_1 _12034_ (.A(_06366_),
    .B(_06365_),
    .Y(_06387_));
 sky130_fd_sc_hd__nor2_1 _12035_ (.A(_06377_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__a32o_1 _12036_ (.A1(_06378_),
    .A2(_06383_),
    .A3(_06384_),
    .B1(_06386_),
    .B2(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__buf_6 _12037_ (.A(\sinegen0.read_ptr[2] ),
    .X(_06390_));
 sky130_fd_sc_hd__buf_2 _12038_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__and3_2 _12039_ (.A(_06391_),
    .B(_06364_),
    .C(_06365_),
    .X(_06392_));
 sky130_fd_sc_hd__o21ai_2 _12040_ (.A1(_06366_),
    .A2(_06364_),
    .B1(_06376_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _12041_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__inv_2 _12042_ (.A(\sinegen0.read_ptr[3] ),
    .Y(_06395_));
 sky130_fd_sc_hd__clkbuf_4 _12043_ (.A(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__clkbuf_4 _12044_ (.A(_06362_),
    .X(_06397_));
 sky130_fd_sc_hd__buf_4 _12045_ (.A(_06366_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_4 _12046_ (.A(_06365_),
    .X(_06399_));
 sky130_fd_sc_hd__nor4_2 _12047_ (.A(_06397_),
    .B(_06398_),
    .C(_06380_),
    .D(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__clkinv_4 _12048_ (.A(\sinegen0.read_ptr[4] ),
    .Y(_06401_));
 sky130_fd_sc_hd__clkbuf_4 _12049_ (.A(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__a211o_1 _12050_ (.A1(_06396_),
    .A2(_06367_),
    .B1(_06400_),
    .C1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_4 _12051_ (.A(\sinegen0.read_ptr[5] ),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_4 _12052_ (.A(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__o221a_1 _12053_ (.A1(_06359_),
    .A2(_06389_),
    .B1(_06394_),
    .B2(_06403_),
    .C1(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__or4_2 _12054_ (.A(_06357_),
    .B(_06371_),
    .C(_06375_),
    .D(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__buf_8 _12055_ (.A(_00004_),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_16 _12056_ (.A(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__buf_12 _12057_ (.A(_00000_),
    .X(_06410_));
 sky130_fd_sc_hd__inv_2 _12058_ (.A(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__buf_4 _12059_ (.A(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__buf_8 _12060_ (.A(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__buf_8 _12061_ (.A(_00000_),
    .X(_06414_));
 sky130_fd_sc_hd__buf_12 _12062_ (.A(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__buf_12 _12063_ (.A(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(_06416_),
    .B(\fifo0.fifo_store[38][15] ),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_16 _12065_ (.A(_00001_),
    .X(_06418_));
 sky130_fd_sc_hd__buf_8 _12066_ (.A(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__buf_12 _12067_ (.A(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__buf_12 _12068_ (.A(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__buf_12 _12069_ (.A(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__o211a_1 _12070_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[39][15] ),
    .B1(_06417_),
    .C1(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__clkinv_8 _12071_ (.A(_06419_),
    .Y(_06424_));
 sky130_fd_sc_hd__buf_12 _12072_ (.A(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_12 _12073_ (.A(_06410_),
    .X(_06426_));
 sky130_fd_sc_hd__buf_6 _12074_ (.A(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__mux2_1 _12075_ (.A0(\fifo0.fifo_store[36][15] ),
    .A1(\fifo0.fifo_store[37][15] ),
    .S(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__inv_2 _12076_ (.A(_00002_),
    .Y(_06429_));
 sky130_fd_sc_hd__buf_6 _12077_ (.A(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__buf_12 _12078_ (.A(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__a21o_1 _12079_ (.A1(_06425_),
    .A2(_06428_),
    .B1(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__buf_8 _12080_ (.A(_06410_),
    .X(_06433_));
 sky130_fd_sc_hd__buf_12 _12081_ (.A(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_12 _12082_ (.A(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__buf_6 _12083_ (.A(_06418_),
    .X(_06436_));
 sky130_fd_sc_hd__buf_12 _12084_ (.A(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__buf_12 _12085_ (.A(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__mux4_1 _12086_ (.A0(\fifo0.fifo_store[32][15] ),
    .A1(\fifo0.fifo_store[33][15] ),
    .A2(\fifo0.fifo_store[34][15] ),
    .A3(\fifo0.fifo_store[35][15] ),
    .S0(_06435_),
    .S1(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_16 _12087_ (.A(_00002_),
    .X(_06440_));
 sky130_fd_sc_hd__buf_12 _12088_ (.A(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_8 _12089_ (.A(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__inv_2 _12090_ (.A(_00003_),
    .Y(_06443_));
 sky130_fd_sc_hd__buf_8 _12091_ (.A(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__buf_8 _12092_ (.A(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__o221a_1 _12093_ (.A1(_06423_),
    .A2(_06432_),
    .B1(_06439_),
    .B2(_06442_),
    .C1(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__buf_12 _12094_ (.A(_00002_),
    .X(_06447_));
 sky130_fd_sc_hd__buf_12 _12095_ (.A(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__buf_12 _12096_ (.A(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__buf_8 _12097_ (.A(_06410_),
    .X(_06450_));
 sky130_fd_sc_hd__buf_12 _12098_ (.A(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__buf_12 _12099_ (.A(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_16 _12100_ (.A(_06436_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_12 _12101_ (.A(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__mux4_1 _12102_ (.A0(\fifo0.fifo_store[40][15] ),
    .A1(\fifo0.fifo_store[41][15] ),
    .A2(\fifo0.fifo_store[42][15] ),
    .A3(\fifo0.fifo_store[43][15] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__buf_8 _12103_ (.A(_06430_),
    .X(_06456_));
 sky130_fd_sc_hd__buf_12 _12104_ (.A(_06433_),
    .X(_06457_));
 sky130_fd_sc_hd__buf_12 _12105_ (.A(_06436_),
    .X(_06458_));
 sky130_fd_sc_hd__mux4_1 _12106_ (.A0(\fifo0.fifo_store[44][15] ),
    .A1(\fifo0.fifo_store[45][15] ),
    .A2(\fifo0.fifo_store[46][15] ),
    .A3(\fifo0.fifo_store[47][15] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__or2_1 _12107_ (.A(_06456_),
    .B(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__buf_8 _12108_ (.A(_00003_),
    .X(_06461_));
 sky130_fd_sc_hd__buf_8 _12109_ (.A(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_16 _12110_ (.A(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__o211a_1 _12111_ (.A1(_06449_),
    .A2(_06455_),
    .B1(_06460_),
    .C1(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__buf_12 _12112_ (.A(_00005_),
    .X(_06465_));
 sky130_fd_sc_hd__clkbuf_16 _12113_ (.A(_06443_),
    .X(_06466_));
 sky130_fd_sc_hd__buf_12 _12114_ (.A(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__buf_8 _12115_ (.A(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__buf_12 _12116_ (.A(_06433_),
    .X(_06469_));
 sky130_fd_sc_hd__buf_6 _12117_ (.A(_06418_),
    .X(_06470_));
 sky130_fd_sc_hd__buf_12 _12118_ (.A(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__mux4_1 _12119_ (.A0(\fifo0.fifo_store[48][15] ),
    .A1(\fifo0.fifo_store[49][15] ),
    .A2(\fifo0.fifo_store[50][15] ),
    .A3(\fifo0.fifo_store[51][15] ),
    .S0(_06469_),
    .S1(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__mux4_1 _12120_ (.A0(\fifo0.fifo_store[52][15] ),
    .A1(\fifo0.fifo_store[53][15] ),
    .A2(\fifo0.fifo_store[54][15] ),
    .A3(\fifo0.fifo_store[55][15] ),
    .S0(_06469_),
    .S1(_06471_),
    .X(_06473_));
 sky130_fd_sc_hd__buf_12 _12121_ (.A(_06440_),
    .X(_06474_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(_06472_),
    .A1(_06473_),
    .S(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_16 _12123_ (.A(_06429_),
    .X(_06476_));
 sky130_fd_sc_hd__buf_8 _12124_ (.A(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__buf_12 _12125_ (.A(_06410_),
    .X(_06478_));
 sky130_fd_sc_hd__buf_12 _12126_ (.A(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__buf_12 _12127_ (.A(_06418_),
    .X(_06480_));
 sky130_fd_sc_hd__buf_12 _12128_ (.A(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__mux4_1 _12129_ (.A0(\fifo0.fifo_store[60][15] ),
    .A1(\fifo0.fifo_store[61][15] ),
    .A2(\fifo0.fifo_store[62][15] ),
    .A3(\fifo0.fifo_store[63][15] ),
    .S0(_06479_),
    .S1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__or2_1 _12130_ (.A(_06477_),
    .B(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__buf_8 _12131_ (.A(_00002_),
    .X(_06484_));
 sky130_fd_sc_hd__clkbuf_16 _12132_ (.A(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__buf_12 _12133_ (.A(_06410_),
    .X(_06486_));
 sky130_fd_sc_hd__buf_12 _12134_ (.A(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__buf_12 _12135_ (.A(_06418_),
    .X(_06488_));
 sky130_fd_sc_hd__buf_12 _12136_ (.A(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__mux4_1 _12137_ (.A0(\fifo0.fifo_store[56][15] ),
    .A1(\fifo0.fifo_store[57][15] ),
    .A2(\fifo0.fifo_store[58][15] ),
    .A3(\fifo0.fifo_store[59][15] ),
    .S0(_06487_),
    .S1(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__buf_6 _12138_ (.A(_06461_),
    .X(_06491_));
 sky130_fd_sc_hd__o21a_1 _12139_ (.A1(_06485_),
    .A2(_06490_),
    .B1(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__inv_8 _12140_ (.A(_00004_),
    .Y(_06493_));
 sky130_fd_sc_hd__buf_12 _12141_ (.A(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__a221o_1 _12142_ (.A1(_06468_),
    .A2(_06475_),
    .B1(_06483_),
    .B2(_06492_),
    .C1(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__o311a_1 _12143_ (.A1(_06409_),
    .A2(_06446_),
    .A3(_06464_),
    .B1(_06465_),
    .C1(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__clkinv_4 _12144_ (.A(_00005_),
    .Y(_06497_));
 sky130_fd_sc_hd__buf_12 _12145_ (.A(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__buf_8 _12146_ (.A(_06433_),
    .X(_06499_));
 sky130_fd_sc_hd__mux4_1 _12147_ (.A0(\fifo0.fifo_store[0][15] ),
    .A1(\fifo0.fifo_store[1][15] ),
    .A2(\fifo0.fifo_store[2][15] ),
    .A3(\fifo0.fifo_store[3][15] ),
    .S0(_06499_),
    .S1(_06437_),
    .X(_06500_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(_06441_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__buf_6 _12149_ (.A(_06430_),
    .X(_06502_));
 sky130_fd_sc_hd__buf_12 _12150_ (.A(_06450_),
    .X(_06503_));
 sky130_fd_sc_hd__buf_12 _12151_ (.A(_06436_),
    .X(_06504_));
 sky130_fd_sc_hd__mux4_1 _12152_ (.A0(\fifo0.fifo_store[4][15] ),
    .A1(\fifo0.fifo_store[5][15] ),
    .A2(\fifo0.fifo_store[6][15] ),
    .A3(\fifo0.fifo_store[7][15] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__o21a_1 _12153_ (.A1(_06502_),
    .A2(_06505_),
    .B1(_06444_),
    .X(_06506_));
 sky130_fd_sc_hd__buf_12 _12154_ (.A(_06414_),
    .X(_06507_));
 sky130_fd_sc_hd__buf_12 _12155_ (.A(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__or2b_1 _12156_ (.A(\fifo0.fifo_store[15][15] ),
    .B_N(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__buf_12 _12157_ (.A(_06418_),
    .X(_06510_));
 sky130_fd_sc_hd__buf_12 _12158_ (.A(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__o21a_1 _12159_ (.A1(_06508_),
    .A2(\fifo0.fifo_store[14][15] ),
    .B1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__buf_12 _12160_ (.A(_06414_),
    .X(_06513_));
 sky130_fd_sc_hd__buf_12 _12161_ (.A(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(\fifo0.fifo_store[12][15] ),
    .A1(\fifo0.fifo_store[13][15] ),
    .S(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__buf_12 _12163_ (.A(_06424_),
    .X(_06516_));
 sky130_fd_sc_hd__buf_8 _12164_ (.A(_06476_),
    .X(_06517_));
 sky130_fd_sc_hd__a221o_1 _12165_ (.A1(_06509_),
    .A2(_06512_),
    .B1(_06515_),
    .B2(_06516_),
    .C1(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__buf_12 _12166_ (.A(_06447_),
    .X(_06519_));
 sky130_fd_sc_hd__buf_12 _12167_ (.A(_06410_),
    .X(_06520_));
 sky130_fd_sc_hd__buf_12 _12168_ (.A(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__buf_8 _12169_ (.A(_06418_),
    .X(_06522_));
 sky130_fd_sc_hd__buf_12 _12170_ (.A(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__mux4_2 _12171_ (.A0(\fifo0.fifo_store[8][15] ),
    .A1(\fifo0.fifo_store[9][15] ),
    .A2(\fifo0.fifo_store[10][15] ),
    .A3(\fifo0.fifo_store[11][15] ),
    .S0(_06521_),
    .S1(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__o21a_1 _12172_ (.A1(_06519_),
    .A2(_06524_),
    .B1(_06462_),
    .X(_06525_));
 sky130_fd_sc_hd__a221o_1 _12173_ (.A1(_06501_),
    .A2(_06506_),
    .B1(_06518_),
    .B2(_06525_),
    .C1(_06408_),
    .X(_06526_));
 sky130_fd_sc_hd__buf_12 _12174_ (.A(_06414_),
    .X(_06527_));
 sky130_fd_sc_hd__buf_12 _12175_ (.A(_06470_),
    .X(_06528_));
 sky130_fd_sc_hd__mux4_1 _12176_ (.A0(\fifo0.fifo_store[16][15] ),
    .A1(\fifo0.fifo_store[17][15] ),
    .A2(\fifo0.fifo_store[18][15] ),
    .A3(\fifo0.fifo_store[19][15] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__mux4_1 _12177_ (.A0(\fifo0.fifo_store[20][15] ),
    .A1(\fifo0.fifo_store[21][15] ),
    .A2(\fifo0.fifo_store[22][15] ),
    .A3(\fifo0.fifo_store[23][15] ),
    .S0(_06507_),
    .S1(_06528_),
    .X(_06530_));
 sky130_fd_sc_hd__clkbuf_16 _12178_ (.A(_06440_),
    .X(_06531_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(_06529_),
    .A1(_06530_),
    .S(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__buf_12 _12180_ (.A(_06450_),
    .X(_06533_));
 sky130_fd_sc_hd__mux4_1 _12181_ (.A0(\fifo0.fifo_store[28][15] ),
    .A1(\fifo0.fifo_store[29][15] ),
    .A2(\fifo0.fifo_store[30][15] ),
    .A3(\fifo0.fifo_store[31][15] ),
    .S0(_06533_),
    .S1(_06458_),
    .X(_06534_));
 sky130_fd_sc_hd__or2_1 _12182_ (.A(_06517_),
    .B(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__buf_12 _12183_ (.A(_06450_),
    .X(_06536_));
 sky130_fd_sc_hd__mux4_1 _12184_ (.A0(\fifo0.fifo_store[24][15] ),
    .A1(\fifo0.fifo_store[25][15] ),
    .A2(\fifo0.fifo_store[26][15] ),
    .A3(\fifo0.fifo_store[27][15] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_06537_));
 sky130_fd_sc_hd__o21a_1 _12185_ (.A1(_06519_),
    .A2(_06537_),
    .B1(_06462_),
    .X(_06538_));
 sky130_fd_sc_hd__buf_12 _12186_ (.A(_06493_),
    .X(_06539_));
 sky130_fd_sc_hd__a221o_1 _12187_ (.A1(_06445_),
    .A2(_06532_),
    .B1(_06535_),
    .B2(_06538_),
    .C1(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__a31o_1 _12188_ (.A1(_06498_),
    .A2(_06526_),
    .A3(_06540_),
    .B1(_00006_),
    .X(_06541_));
 sky130_fd_sc_hd__buf_12 _12189_ (.A(_06469_),
    .X(_06542_));
 sky130_fd_sc_hd__mux4_2 _12190_ (.A0(\fifo0.fifo_store[96][15] ),
    .A1(\fifo0.fifo_store[97][15] ),
    .A2(\fifo0.fifo_store[98][15] ),
    .A3(\fifo0.fifo_store[99][15] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_06543_));
 sky130_fd_sc_hd__buf_12 _12191_ (.A(_06414_),
    .X(_06544_));
 sky130_fd_sc_hd__clkbuf_16 _12192_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__or2b_1 _12193_ (.A(\fifo0.fifo_store[103][15] ),
    .B_N(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__o21a_1 _12194_ (.A1(_06545_),
    .A2(\fifo0.fifo_store[102][15] ),
    .B1(_06489_),
    .X(_06547_));
 sky130_fd_sc_hd__buf_12 _12195_ (.A(_06410_),
    .X(_06548_));
 sky130_fd_sc_hd__clkbuf_16 _12196_ (.A(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(\fifo0.fifo_store[100][15] ),
    .A1(\fifo0.fifo_store[101][15] ),
    .S(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__a221o_1 _12198_ (.A1(_06546_),
    .A2(_06547_),
    .B1(_06550_),
    .B2(_06516_),
    .C1(_06431_),
    .X(_06551_));
 sky130_fd_sc_hd__buf_12 _12199_ (.A(_06467_),
    .X(_06552_));
 sky130_fd_sc_hd__o211a_1 _12200_ (.A1(_06449_),
    .A2(_06543_),
    .B1(_06551_),
    .C1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__buf_8 _12201_ (.A(_06448_),
    .X(_06554_));
 sky130_fd_sc_hd__buf_12 _12202_ (.A(_06522_),
    .X(_06555_));
 sky130_fd_sc_hd__buf_12 _12203_ (.A(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__mux4_1 _12204_ (.A0(\fifo0.fifo_store[104][15] ),
    .A1(\fifo0.fifo_store[105][15] ),
    .A2(\fifo0.fifo_store[106][15] ),
    .A3(\fifo0.fifo_store[107][15] ),
    .S0(_06452_),
    .S1(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__mux4_1 _12205_ (.A0(\fifo0.fifo_store[108][15] ),
    .A1(\fifo0.fifo_store[109][15] ),
    .A2(\fifo0.fifo_store[110][15] ),
    .A3(\fifo0.fifo_store[111][15] ),
    .S0(_06457_),
    .S1(_06453_),
    .X(_06558_));
 sky130_fd_sc_hd__or2_1 _12206_ (.A(_06456_),
    .B(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__o211a_1 _12207_ (.A1(_06554_),
    .A2(_06557_),
    .B1(_06559_),
    .C1(_06463_),
    .X(_06560_));
 sky130_fd_sc_hd__buf_12 _12208_ (.A(_06470_),
    .X(_06561_));
 sky130_fd_sc_hd__mux4_1 _12209_ (.A0(\fifo0.fifo_store[112][15] ),
    .A1(\fifo0.fifo_store[113][15] ),
    .A2(\fifo0.fifo_store[114][15] ),
    .A3(\fifo0.fifo_store[115][15] ),
    .S0(_06434_),
    .S1(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__buf_12 _12210_ (.A(_06433_),
    .X(_06563_));
 sky130_fd_sc_hd__mux4_1 _12211_ (.A0(\fifo0.fifo_store[116][15] ),
    .A1(\fifo0.fifo_store[117][15] ),
    .A2(\fifo0.fifo_store[118][15] ),
    .A3(\fifo0.fifo_store[119][15] ),
    .S0(_06563_),
    .S1(_06561_),
    .X(_06564_));
 sky130_fd_sc_hd__buf_12 _12212_ (.A(_06440_),
    .X(_06565_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(_06562_),
    .A1(_06564_),
    .S(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__mux4_1 _12214_ (.A0(\fifo0.fifo_store[124][15] ),
    .A1(\fifo0.fifo_store[125][15] ),
    .A2(\fifo0.fifo_store[126][15] ),
    .A3(\fifo0.fifo_store[127][15] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_06567_));
 sky130_fd_sc_hd__or2_1 _12215_ (.A(_06502_),
    .B(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__buf_12 _12216_ (.A(_06520_),
    .X(_06569_));
 sky130_fd_sc_hd__mux4_2 _12217_ (.A0(\fifo0.fifo_store[120][15] ),
    .A1(\fifo0.fifo_store[121][15] ),
    .A2(\fifo0.fifo_store[122][15] ),
    .A3(\fifo0.fifo_store[123][15] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_06570_));
 sky130_fd_sc_hd__buf_12 _12218_ (.A(_06461_),
    .X(_06571_));
 sky130_fd_sc_hd__o21a_1 _12219_ (.A1(_06485_),
    .A2(_06570_),
    .B1(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__a221o_1 _12220_ (.A1(_06552_),
    .A2(_06566_),
    .B1(_06568_),
    .B2(_06572_),
    .C1(_06494_),
    .X(_06573_));
 sky130_fd_sc_hd__o311a_4 _12221_ (.A1(_06409_),
    .A2(_06553_),
    .A3(_06560_),
    .B1(_06573_),
    .C1(_06465_),
    .X(_06574_));
 sky130_fd_sc_hd__buf_12 _12222_ (.A(_06497_),
    .X(_06575_));
 sky130_fd_sc_hd__buf_12 _12223_ (.A(_06544_),
    .X(_06576_));
 sky130_fd_sc_hd__or2b_1 _12224_ (.A(\fifo0.fifo_store[79][15] ),
    .B_N(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__buf_12 _12225_ (.A(_06418_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_12 _12226_ (.A(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__o21a_1 _12227_ (.A1(_06576_),
    .A2(\fifo0.fifo_store[78][15] ),
    .B1(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _12228_ (.A0(\fifo0.fifo_store[76][15] ),
    .A1(\fifo0.fifo_store[77][15] ),
    .S(_06514_),
    .X(_06581_));
 sky130_fd_sc_hd__a221o_1 _12229_ (.A1(_06577_),
    .A2(_06580_),
    .B1(_06581_),
    .B2(_06516_),
    .C1(_06517_),
    .X(_06582_));
 sky130_fd_sc_hd__mux4_1 _12230_ (.A0(\fifo0.fifo_store[72][15] ),
    .A1(\fifo0.fifo_store[73][15] ),
    .A2(\fifo0.fifo_store[74][15] ),
    .A3(\fifo0.fifo_store[75][15] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_06583_));
 sky130_fd_sc_hd__o21a_1 _12231_ (.A1(_06519_),
    .A2(_06583_),
    .B1(_06462_),
    .X(_06584_));
 sky130_fd_sc_hd__mux4_2 _12232_ (.A0(\fifo0.fifo_store[64][15] ),
    .A1(\fifo0.fifo_store[65][15] ),
    .A2(\fifo0.fifo_store[66][15] ),
    .A3(\fifo0.fifo_store[67][15] ),
    .S0(_06469_),
    .S1(_06471_),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_16 _12233_ (.A(_06433_),
    .X(_06586_));
 sky130_fd_sc_hd__mux4_1 _12234_ (.A0(\fifo0.fifo_store[68][15] ),
    .A1(\fifo0.fifo_store[69][15] ),
    .A2(\fifo0.fifo_store[70][15] ),
    .A3(\fifo0.fifo_store[71][15] ),
    .S0(_06586_),
    .S1(_06471_),
    .X(_06587_));
 sky130_fd_sc_hd__mux2_2 _12235_ (.A0(_06585_),
    .A1(_06587_),
    .S(_06474_),
    .X(_06588_));
 sky130_fd_sc_hd__buf_8 _12236_ (.A(_00004_),
    .X(_06589_));
 sky130_fd_sc_hd__a221o_1 _12237_ (.A1(_06582_),
    .A2(_06584_),
    .B1(_06588_),
    .B2(_06445_),
    .C1(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__buf_12 _12238_ (.A(_06433_),
    .X(_06591_));
 sky130_fd_sc_hd__buf_8 _12239_ (.A(_06436_),
    .X(_06592_));
 sky130_fd_sc_hd__mux4_1 _12240_ (.A0(\fifo0.fifo_store[88][15] ),
    .A1(\fifo0.fifo_store[89][15] ),
    .A2(\fifo0.fifo_store[90][15] ),
    .A3(\fifo0.fifo_store[91][15] ),
    .S0(_06591_),
    .S1(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__or2_1 _12241_ (.A(_06448_),
    .B(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__mux4_2 _12242_ (.A0(\fifo0.fifo_store[92][15] ),
    .A1(\fifo0.fifo_store[93][15] ),
    .A2(\fifo0.fifo_store[94][15] ),
    .A3(\fifo0.fifo_store[95][15] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_06595_));
 sky130_fd_sc_hd__o21a_1 _12243_ (.A1(_06477_),
    .A2(_06595_),
    .B1(_06462_),
    .X(_06596_));
 sky130_fd_sc_hd__mux4_1 _12244_ (.A0(\fifo0.fifo_store[84][15] ),
    .A1(\fifo0.fifo_store[85][15] ),
    .A2(\fifo0.fifo_store[86][15] ),
    .A3(\fifo0.fifo_store[87][15] ),
    .S0(_06451_),
    .S1(_06453_),
    .X(_06597_));
 sky130_fd_sc_hd__or2_1 _12245_ (.A(_06456_),
    .B(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__buf_12 _12246_ (.A(_06484_),
    .X(_06599_));
 sky130_fd_sc_hd__buf_12 _12247_ (.A(_06520_),
    .X(_06600_));
 sky130_fd_sc_hd__mux4_1 _12248_ (.A0(\fifo0.fifo_store[80][15] ),
    .A1(\fifo0.fifo_store[81][15] ),
    .A2(\fifo0.fifo_store[82][15] ),
    .A3(\fifo0.fifo_store[83][15] ),
    .S0(_06600_),
    .S1(_06555_),
    .X(_06601_));
 sky130_fd_sc_hd__o21a_1 _12249_ (.A1(_06599_),
    .A2(_06601_),
    .B1(_06467_),
    .X(_06602_));
 sky130_fd_sc_hd__a221o_1 _12250_ (.A1(_06594_),
    .A2(_06596_),
    .B1(_06598_),
    .B2(_06602_),
    .C1(_06539_),
    .X(_06603_));
 sky130_fd_sc_hd__clkinv_8 _12251_ (.A(_00006_),
    .Y(_06604_));
 sky130_fd_sc_hd__a31o_2 _12252_ (.A1(_06575_),
    .A2(_06590_),
    .A3(_06603_),
    .B1(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__buf_6 _12253_ (.A(_06357_),
    .X(_06606_));
 sky130_fd_sc_hd__o221ai_4 _12254_ (.A1(_06496_),
    .A2(_06541_),
    .B1(_06574_),
    .B2(_06605_),
    .C1(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__and2_1 _12255_ (.A(_06407_),
    .B(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__nor2_2 _12256_ (.A(_06356_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__xnor2_1 _12257_ (.A(\dsmod0.accu1[15] ),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__buf_4 _12258_ (.A(_06357_),
    .X(_06611_));
 sky130_fd_sc_hd__buf_8 _12259_ (.A(_06411_),
    .X(_06612_));
 sky130_fd_sc_hd__or2_1 _12260_ (.A(_06544_),
    .B(\fifo0.fifo_store[54][14] ),
    .X(_06613_));
 sky130_fd_sc_hd__buf_12 _12261_ (.A(_06419_),
    .X(_06614_));
 sky130_fd_sc_hd__buf_12 _12262_ (.A(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__o211a_1 _12263_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[55][14] ),
    .B1(_06613_),
    .C1(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_12 _12264_ (.A(_06414_),
    .X(_06617_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(\fifo0.fifo_store[52][14] ),
    .A1(\fifo0.fifo_store[53][14] ),
    .S(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(_06424_),
    .A2(_06618_),
    .B1(_06476_),
    .X(_06619_));
 sky130_fd_sc_hd__mux4_1 _12267_ (.A0(\fifo0.fifo_store[48][14] ),
    .A1(\fifo0.fifo_store[49][14] ),
    .A2(\fifo0.fifo_store[50][14] ),
    .A3(\fifo0.fifo_store[51][14] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_06620_));
 sky130_fd_sc_hd__buf_8 _12268_ (.A(_06466_),
    .X(_06621_));
 sky130_fd_sc_hd__o221a_1 _12269_ (.A1(_06616_),
    .A2(_06619_),
    .B1(_06620_),
    .B2(_06519_),
    .C1(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__buf_8 _12270_ (.A(_00002_),
    .X(_06623_));
 sky130_fd_sc_hd__buf_12 _12271_ (.A(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__buf_12 _12272_ (.A(_06486_),
    .X(_06625_));
 sky130_fd_sc_hd__mux4_1 _12273_ (.A0(\fifo0.fifo_store[56][14] ),
    .A1(\fifo0.fifo_store[57][14] ),
    .A2(\fifo0.fifo_store[58][14] ),
    .A3(\fifo0.fifo_store[59][14] ),
    .S0(_06625_),
    .S1(_06489_),
    .X(_06626_));
 sky130_fd_sc_hd__buf_12 _12274_ (.A(_06418_),
    .X(_06627_));
 sky130_fd_sc_hd__mux4_1 _12275_ (.A0(\fifo0.fifo_store[60][14] ),
    .A1(\fifo0.fifo_store[61][14] ),
    .A2(\fifo0.fifo_store[62][14] ),
    .A3(\fifo0.fifo_store[63][14] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__or2_1 _12276_ (.A(_06476_),
    .B(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__buf_8 _12277_ (.A(_06461_),
    .X(_06630_));
 sky130_fd_sc_hd__o211a_1 _12278_ (.A1(_06624_),
    .A2(_06626_),
    .B1(_06629_),
    .C1(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__mux4_1 _12279_ (.A0(\fifo0.fifo_store[40][14] ),
    .A1(\fifo0.fifo_store[41][14] ),
    .A2(\fifo0.fifo_store[42][14] ),
    .A3(\fifo0.fifo_store[43][14] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_06632_));
 sky130_fd_sc_hd__or2_1 _12280_ (.A(_06484_),
    .B(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__buf_8 _12281_ (.A(_06429_),
    .X(_06634_));
 sky130_fd_sc_hd__mux4_2 _12282_ (.A0(\fifo0.fifo_store[44][14] ),
    .A1(\fifo0.fifo_store[45][14] ),
    .A2(\fifo0.fifo_store[46][14] ),
    .A3(\fifo0.fifo_store[47][14] ),
    .S0(_06426_),
    .S1(_06488_),
    .X(_06635_));
 sky130_fd_sc_hd__o21a_1 _12283_ (.A1(_06634_),
    .A2(_06635_),
    .B1(_06461_),
    .X(_06636_));
 sky130_fd_sc_hd__mux4_2 _12284_ (.A0(\fifo0.fifo_store[32][14] ),
    .A1(\fifo0.fifo_store[33][14] ),
    .A2(\fifo0.fifo_store[34][14] ),
    .A3(\fifo0.fifo_store[35][14] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_06637_));
 sky130_fd_sc_hd__or2_1 _12285_ (.A(_06484_),
    .B(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__mux4_1 _12286_ (.A0(\fifo0.fifo_store[36][14] ),
    .A1(\fifo0.fifo_store[37][14] ),
    .A2(\fifo0.fifo_store[38][14] ),
    .A3(\fifo0.fifo_store[39][14] ),
    .S0(_06426_),
    .S1(_06578_),
    .X(_06639_));
 sky130_fd_sc_hd__o21a_1 _12287_ (.A1(_06634_),
    .A2(_06639_),
    .B1(_06466_),
    .X(_06640_));
 sky130_fd_sc_hd__buf_12 _12288_ (.A(_00004_),
    .X(_06641_));
 sky130_fd_sc_hd__a221o_1 _12289_ (.A1(_06633_),
    .A2(_06636_),
    .B1(_06638_),
    .B2(_06640_),
    .C1(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__buf_12 _12290_ (.A(_00005_),
    .X(_06643_));
 sky130_fd_sc_hd__o311a_1 _12291_ (.A1(_06494_),
    .A2(_06622_),
    .A3(_06631_),
    .B1(_06642_),
    .C1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__buf_12 _12292_ (.A(_06433_),
    .X(_06645_));
 sky130_fd_sc_hd__or2_1 _12293_ (.A(_06645_),
    .B(\fifo0.fifo_store[6][14] ),
    .X(_06646_));
 sky130_fd_sc_hd__clkbuf_16 _12294_ (.A(_06419_),
    .X(_06647_));
 sky130_fd_sc_hd__buf_12 _12295_ (.A(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__o211a_1 _12296_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[7][14] ),
    .B1(_06646_),
    .C1(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__buf_6 _12297_ (.A(_06424_),
    .X(_06650_));
 sky130_fd_sc_hd__mux2_1 _12298_ (.A0(\fifo0.fifo_store[4][14] ),
    .A1(\fifo0.fifo_store[5][14] ),
    .S(_06415_),
    .X(_06651_));
 sky130_fd_sc_hd__a21o_1 _12299_ (.A1(_06650_),
    .A2(_06651_),
    .B1(_06476_),
    .X(_06652_));
 sky130_fd_sc_hd__mux4_1 _12300_ (.A0(\fifo0.fifo_store[0][14] ),
    .A1(\fifo0.fifo_store[1][14] ),
    .A2(\fifo0.fifo_store[2][14] ),
    .A3(\fifo0.fifo_store[3][14] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_06653_));
 sky130_fd_sc_hd__o221a_1 _12301_ (.A1(_06649_),
    .A2(_06652_),
    .B1(_06653_),
    .B2(_06485_),
    .C1(_06621_),
    .X(_06654_));
 sky130_fd_sc_hd__buf_8 _12302_ (.A(_00002_),
    .X(_06655_));
 sky130_fd_sc_hd__buf_8 _12303_ (.A(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__buf_12 _12304_ (.A(_06410_),
    .X(_06657_));
 sky130_fd_sc_hd__buf_12 _12305_ (.A(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__mux4_2 _12306_ (.A0(\fifo0.fifo_store[8][14] ),
    .A1(\fifo0.fifo_store[9][14] ),
    .A2(\fifo0.fifo_store[10][14] ),
    .A3(\fifo0.fifo_store[11][14] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_06659_));
 sky130_fd_sc_hd__clkbuf_16 _12307_ (.A(_06429_),
    .X(_06660_));
 sky130_fd_sc_hd__mux4_2 _12308_ (.A0(\fifo0.fifo_store[12][14] ),
    .A1(\fifo0.fifo_store[13][14] ),
    .A2(\fifo0.fifo_store[14][14] ),
    .A3(\fifo0.fifo_store[15][14] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_06661_));
 sky130_fd_sc_hd__or2_1 _12309_ (.A(_06660_),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_16 _12310_ (.A(_00003_),
    .X(_06663_));
 sky130_fd_sc_hd__buf_8 _12311_ (.A(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__o211a_1 _12312_ (.A1(_06656_),
    .A2(_06659_),
    .B1(_06662_),
    .C1(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__mux4_1 _12313_ (.A0(\fifo0.fifo_store[24][14] ),
    .A1(\fifo0.fifo_store[25][14] ),
    .A2(\fifo0.fifo_store[26][14] ),
    .A3(\fifo0.fifo_store[27][14] ),
    .S0(_06426_),
    .S1(_06488_),
    .X(_06666_));
 sky130_fd_sc_hd__or2_1 _12314_ (.A(_06623_),
    .B(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__buf_8 _12315_ (.A(_06429_),
    .X(_06668_));
 sky130_fd_sc_hd__mux4_1 _12316_ (.A0(\fifo0.fifo_store[28][14] ),
    .A1(\fifo0.fifo_store[29][14] ),
    .A2(\fifo0.fifo_store[30][14] ),
    .A3(\fifo0.fifo_store[31][14] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_06669_));
 sky130_fd_sc_hd__o21a_1 _12317_ (.A1(_06668_),
    .A2(_06669_),
    .B1(_06461_),
    .X(_06670_));
 sky130_fd_sc_hd__mux4_1 _12318_ (.A0(\fifo0.fifo_store[16][14] ),
    .A1(\fifo0.fifo_store[17][14] ),
    .A2(\fifo0.fifo_store[18][14] ),
    .A3(\fifo0.fifo_store[19][14] ),
    .S0(_06426_),
    .S1(_06578_),
    .X(_06671_));
 sky130_fd_sc_hd__or2_1 _12319_ (.A(_06623_),
    .B(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__buf_12 _12320_ (.A(_06410_),
    .X(_06673_));
 sky130_fd_sc_hd__mux4_1 _12321_ (.A0(\fifo0.fifo_store[20][14] ),
    .A1(\fifo0.fifo_store[21][14] ),
    .A2(\fifo0.fifo_store[22][14] ),
    .A3(\fifo0.fifo_store[23][14] ),
    .S0(_06673_),
    .S1(_06420_),
    .X(_06674_));
 sky130_fd_sc_hd__o21a_1 _12322_ (.A1(_06668_),
    .A2(_06674_),
    .B1(_06466_),
    .X(_06675_));
 sky130_fd_sc_hd__a221o_1 _12323_ (.A1(_06667_),
    .A2(_06670_),
    .B1(_06672_),
    .B2(_06675_),
    .C1(_06493_),
    .X(_06676_));
 sky130_fd_sc_hd__clkbuf_16 _12324_ (.A(_06497_),
    .X(_06677_));
 sky130_fd_sc_hd__o311a_1 _12325_ (.A1(_06589_),
    .A2(_06654_),
    .A3(_06665_),
    .B1(_06676_),
    .C1(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__buf_8 _12326_ (.A(_06493_),
    .X(_06679_));
 sky130_fd_sc_hd__buf_6 _12327_ (.A(_06430_),
    .X(_06680_));
 sky130_fd_sc_hd__buf_6 _12328_ (.A(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__mux4_1 _12329_ (.A0(\fifo0.fifo_store[124][14] ),
    .A1(\fifo0.fifo_store[125][14] ),
    .A2(\fifo0.fifo_store[126][14] ),
    .A3(\fifo0.fifo_store[127][14] ),
    .S0(_06514_),
    .S1(_06615_),
    .X(_06682_));
 sky130_fd_sc_hd__buf_8 _12330_ (.A(_06440_),
    .X(_06683_));
 sky130_fd_sc_hd__mux4_1 _12331_ (.A0(\fifo0.fifo_store[120][14] ),
    .A1(\fifo0.fifo_store[121][14] ),
    .A2(\fifo0.fifo_store[122][14] ),
    .A3(\fifo0.fifo_store[123][14] ),
    .S0(_06548_),
    .S1(_06614_),
    .X(_06684_));
 sky130_fd_sc_hd__or2_1 _12332_ (.A(_06683_),
    .B(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__buf_8 _12333_ (.A(_06663_),
    .X(_06686_));
 sky130_fd_sc_hd__o211a_1 _12334_ (.A1(_06681_),
    .A2(_06682_),
    .B1(_06685_),
    .C1(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__buf_8 _12335_ (.A(_06531_),
    .X(_06688_));
 sky130_fd_sc_hd__buf_12 _12336_ (.A(_06617_),
    .X(_06689_));
 sky130_fd_sc_hd__buf_12 _12337_ (.A(_06419_),
    .X(_06690_));
 sky130_fd_sc_hd__buf_12 _12338_ (.A(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__mux4_1 _12339_ (.A0(\fifo0.fifo_store[112][14] ),
    .A1(\fifo0.fifo_store[113][14] ),
    .A2(\fifo0.fifo_store[114][14] ),
    .A3(\fifo0.fifo_store[115][14] ),
    .S0(_06689_),
    .S1(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__buf_12 _12340_ (.A(_06426_),
    .X(_06693_));
 sky130_fd_sc_hd__or2b_1 _12341_ (.A(\fifo0.fifo_store[119][14] ),
    .B_N(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__buf_12 _12342_ (.A(_06470_),
    .X(_06695_));
 sky130_fd_sc_hd__o21a_1 _12343_ (.A1(_06693_),
    .A2(\fifo0.fifo_store[118][14] ),
    .B1(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__buf_12 _12344_ (.A(_06433_),
    .X(_06697_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(\fifo0.fifo_store[116][14] ),
    .A1(\fifo0.fifo_store[117][14] ),
    .S(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__buf_8 _12346_ (.A(_06424_),
    .X(_06699_));
 sky130_fd_sc_hd__a221o_1 _12347_ (.A1(_06694_),
    .A2(_06696_),
    .B1(_06698_),
    .B2(_06699_),
    .C1(_06680_),
    .X(_06700_));
 sky130_fd_sc_hd__buf_8 _12348_ (.A(_06444_),
    .X(_06701_));
 sky130_fd_sc_hd__o211a_1 _12349_ (.A1(_06688_),
    .A2(_06692_),
    .B1(_06700_),
    .C1(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_16 _12350_ (.A(_06419_),
    .X(_06703_));
 sky130_fd_sc_hd__mux4_2 _12351_ (.A0(\fifo0.fifo_store[96][14] ),
    .A1(\fifo0.fifo_store[97][14] ),
    .A2(\fifo0.fifo_store[98][14] ),
    .A3(\fifo0.fifo_store[99][14] ),
    .S0(_06548_),
    .S1(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__mux4_1 _12352_ (.A0(\fifo0.fifo_store[100][14] ),
    .A1(\fifo0.fifo_store[101][14] ),
    .A2(\fifo0.fifo_store[102][14] ),
    .A3(\fifo0.fifo_store[103][14] ),
    .S0(_06548_),
    .S1(_06614_),
    .X(_06705_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(_06704_),
    .A1(_06705_),
    .S(_06484_),
    .X(_06706_));
 sky130_fd_sc_hd__mux4_1 _12354_ (.A0(\fifo0.fifo_store[104][14] ),
    .A1(\fifo0.fifo_store[105][14] ),
    .A2(\fifo0.fifo_store[106][14] ),
    .A3(\fifo0.fifo_store[107][14] ),
    .S0(_06617_),
    .S1(_06690_),
    .X(_06707_));
 sky130_fd_sc_hd__or2_1 _12355_ (.A(_06531_),
    .B(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__buf_8 _12356_ (.A(_06430_),
    .X(_06709_));
 sky130_fd_sc_hd__buf_12 _12357_ (.A(_06414_),
    .X(_06710_));
 sky130_fd_sc_hd__buf_12 _12358_ (.A(_06419_),
    .X(_06711_));
 sky130_fd_sc_hd__mux4_2 _12359_ (.A0(\fifo0.fifo_store[108][14] ),
    .A1(\fifo0.fifo_store[109][14] ),
    .A2(\fifo0.fifo_store[110][14] ),
    .A3(\fifo0.fifo_store[111][14] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__buf_8 _12360_ (.A(_06461_),
    .X(_06713_));
 sky130_fd_sc_hd__o21a_1 _12361_ (.A1(_06709_),
    .A2(_06712_),
    .B1(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__a221o_1 _12362_ (.A1(_06701_),
    .A2(_06706_),
    .B1(_06708_),
    .B2(_06714_),
    .C1(_06408_),
    .X(_06715_));
 sky130_fd_sc_hd__o311a_2 _12363_ (.A1(_06679_),
    .A2(_06687_),
    .A3(_06702_),
    .B1(_06643_),
    .C1(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__buf_12 _12364_ (.A(_06414_),
    .X(_06717_));
 sky130_fd_sc_hd__buf_12 _12365_ (.A(_06419_),
    .X(_06718_));
 sky130_fd_sc_hd__mux4_1 _12366_ (.A0(\fifo0.fifo_store[72][14] ),
    .A1(\fifo0.fifo_store[73][14] ),
    .A2(\fifo0.fifo_store[74][14] ),
    .A3(\fifo0.fifo_store[75][14] ),
    .S0(_06717_),
    .S1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__or2_1 _12367_ (.A(_06683_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__buf_8 _12368_ (.A(_06430_),
    .X(_06721_));
 sky130_fd_sc_hd__mux4_1 _12369_ (.A0(\fifo0.fifo_store[76][14] ),
    .A1(\fifo0.fifo_store[77][14] ),
    .A2(\fifo0.fifo_store[78][14] ),
    .A3(\fifo0.fifo_store[79][14] ),
    .S0(_06513_),
    .S1(_06647_),
    .X(_06722_));
 sky130_fd_sc_hd__o21a_1 _12370_ (.A1(_06721_),
    .A2(_06722_),
    .B1(_06663_),
    .X(_06723_));
 sky130_fd_sc_hd__or2b_1 _12371_ (.A(\fifo0.fifo_store[71][14] ),
    .B_N(_06625_),
    .X(_06724_));
 sky130_fd_sc_hd__buf_12 _12372_ (.A(_06470_),
    .X(_06725_));
 sky130_fd_sc_hd__o21a_1 _12373_ (.A1(_06625_),
    .A2(\fifo0.fifo_store[70][14] ),
    .B1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(\fifo0.fifo_store[68][14] ),
    .A1(\fifo0.fifo_store[69][14] ),
    .S(_06434_),
    .X(_06727_));
 sky130_fd_sc_hd__buf_6 _12375_ (.A(_06424_),
    .X(_06728_));
 sky130_fd_sc_hd__a221o_1 _12376_ (.A1(_06724_),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06728_),
    .C1(_06680_),
    .X(_06729_));
 sky130_fd_sc_hd__buf_8 _12377_ (.A(_06440_),
    .X(_06730_));
 sky130_fd_sc_hd__buf_12 _12378_ (.A(_06419_),
    .X(_06731_));
 sky130_fd_sc_hd__mux4_2 _12379_ (.A0(\fifo0.fifo_store[64][14] ),
    .A1(\fifo0.fifo_store[65][14] ),
    .A2(\fifo0.fifo_store[66][14] ),
    .A3(\fifo0.fifo_store[67][14] ),
    .S0(_06617_),
    .S1(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__o21a_1 _12380_ (.A1(_06730_),
    .A2(_06732_),
    .B1(_06444_),
    .X(_06733_));
 sky130_fd_sc_hd__a221o_1 _12381_ (.A1(_06720_),
    .A2(_06723_),
    .B1(_06729_),
    .B2(_06733_),
    .C1(_06641_),
    .X(_06734_));
 sky130_fd_sc_hd__buf_8 _12382_ (.A(_06466_),
    .X(_06735_));
 sky130_fd_sc_hd__mux4_1 _12383_ (.A0(\fifo0.fifo_store[80][14] ),
    .A1(\fifo0.fifo_store[81][14] ),
    .A2(\fifo0.fifo_store[82][14] ),
    .A3(\fifo0.fifo_store[83][14] ),
    .S0(_06426_),
    .S1(_06578_),
    .X(_06736_));
 sky130_fd_sc_hd__mux4_1 _12384_ (.A0(\fifo0.fifo_store[84][14] ),
    .A1(\fifo0.fifo_store[85][14] ),
    .A2(\fifo0.fifo_store[86][14] ),
    .A3(\fifo0.fifo_store[87][14] ),
    .S0(_06426_),
    .S1(_06488_),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(_06736_),
    .A1(_06737_),
    .S(_06447_),
    .X(_06738_));
 sky130_fd_sc_hd__mux4_1 _12386_ (.A0(\fifo0.fifo_store[88][14] ),
    .A1(\fifo0.fifo_store[89][14] ),
    .A2(\fifo0.fifo_store[90][14] ),
    .A3(\fifo0.fifo_store[91][14] ),
    .S0(_06513_),
    .S1(_06718_),
    .X(_06739_));
 sky130_fd_sc_hd__or2_1 _12387_ (.A(_06730_),
    .B(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__mux4_1 _12388_ (.A0(\fifo0.fifo_store[92][14] ),
    .A1(\fifo0.fifo_store[93][14] ),
    .A2(\fifo0.fifo_store[94][14] ),
    .A3(\fifo0.fifo_store[95][14] ),
    .S0(_06513_),
    .S1(_06731_),
    .X(_06741_));
 sky130_fd_sc_hd__o21a_1 _12389_ (.A1(_06721_),
    .A2(_06741_),
    .B1(_06663_),
    .X(_06742_));
 sky130_fd_sc_hd__buf_6 _12390_ (.A(_06493_),
    .X(_06743_));
 sky130_fd_sc_hd__a221o_2 _12391_ (.A1(_06735_),
    .A2(_06738_),
    .B1(_06740_),
    .B2(_06742_),
    .C1(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__a31o_1 _12392_ (.A1(_06677_),
    .A2(_06734_),
    .A3(_06744_),
    .B1(_06604_),
    .X(_06745_));
 sky130_fd_sc_hd__o32a_4 _12393_ (.A1(_00006_),
    .A2(_06644_),
    .A3(_06678_),
    .B1(_06716_),
    .B2(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__buf_2 _12394_ (.A(\sinegen0.read_ptr[6] ),
    .X(_06747_));
 sky130_fd_sc_hd__clkinv_4 _12395_ (.A(_06390_),
    .Y(_06748_));
 sky130_fd_sc_hd__a211o_1 _12396_ (.A1(_06748_),
    .A2(_06361_),
    .B1(_06382_),
    .C1(_06377_),
    .X(_06749_));
 sky130_fd_sc_hd__xor2_1 _12397_ (.A(\sinegen0.read_ptr[1] ),
    .B(\sinegen0.read_ptr[0] ),
    .X(_06750_));
 sky130_fd_sc_hd__clkbuf_4 _12398_ (.A(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__a21o_1 _12399_ (.A1(_06748_),
    .A2(_06751_),
    .B1(_06395_),
    .X(_06752_));
 sky130_fd_sc_hd__nand2_4 _12400_ (.A(\sinegen0.read_ptr[2] ),
    .B(\sinegen0.read_ptr[1] ),
    .Y(_06753_));
 sky130_fd_sc_hd__or2_1 _12401_ (.A(_06377_),
    .B(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__a31o_1 _12402_ (.A1(_06749_),
    .A2(_06752_),
    .A3(_06754_),
    .B1(_06402_),
    .X(_06755_));
 sky130_fd_sc_hd__buf_4 _12403_ (.A(\sinegen0.read_ptr[0] ),
    .X(_06756_));
 sky130_fd_sc_hd__or3_2 _12404_ (.A(_06390_),
    .B(_06379_),
    .C(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__nor2_1 _12405_ (.A(_06396_),
    .B(_06367_),
    .Y(_06758_));
 sky130_fd_sc_hd__and2b_2 _12406_ (.A_N(_06379_),
    .B(_06756_),
    .X(_06759_));
 sky130_fd_sc_hd__a21o_1 _12407_ (.A1(_06395_),
    .A2(_06759_),
    .B1(_06373_),
    .X(_06760_));
 sky130_fd_sc_hd__nand2b_2 _12408_ (.A_N(_06756_),
    .B(_06379_),
    .Y(_06761_));
 sky130_fd_sc_hd__a21oi_2 _12409_ (.A1(_06398_),
    .A2(_06761_),
    .B1(_06397_),
    .Y(_06762_));
 sky130_fd_sc_hd__a211o_1 _12410_ (.A1(_06757_),
    .A2(_06758_),
    .B1(_06760_),
    .C1(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__nand2_1 _12411_ (.A(_06377_),
    .B(_06380_),
    .Y(_06764_));
 sky130_fd_sc_hd__or2b_1 _12412_ (.A(\sinegen0.read_ptr[0] ),
    .B_N(\sinegen0.read_ptr[2] ),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_4 _12413_ (.A(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__a21o_1 _12414_ (.A1(_06764_),
    .A2(_06766_),
    .B1(_06373_),
    .X(_06767_));
 sky130_fd_sc_hd__or3b_2 _12415_ (.A(_06362_),
    .B(_06364_),
    .C_N(_06391_),
    .X(_06768_));
 sky130_fd_sc_hd__inv_2 _12416_ (.A(\sinegen0.read_ptr[6] ),
    .Y(_06769_));
 sky130_fd_sc_hd__o2111a_1 _12417_ (.A1(_06398_),
    .A2(_06361_),
    .B1(_06767_),
    .C1(_06768_),
    .D1(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__a31o_1 _12418_ (.A1(_06747_),
    .A2(_06755_),
    .A3(_06763_),
    .B1(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__or3_1 _12419_ (.A(_06395_),
    .B(_06391_),
    .C(_06750_),
    .X(_06772_));
 sky130_fd_sc_hd__o311a_1 _12420_ (.A1(_06362_),
    .A2(_06380_),
    .A3(_06382_),
    .B1(_06372_),
    .C1(_06373_),
    .X(_06773_));
 sky130_fd_sc_hd__nor2_1 _12421_ (.A(_06364_),
    .B(_06365_),
    .Y(_06774_));
 sky130_fd_sc_hd__nand2_2 _12422_ (.A(_06376_),
    .B(_06366_),
    .Y(_06775_));
 sky130_fd_sc_hd__o22ai_1 _12423_ (.A1(_06382_),
    .A2(_06774_),
    .B1(_06775_),
    .B2(_06399_),
    .Y(_06776_));
 sky130_fd_sc_hd__o2bb2a_1 _12424_ (.A1_N(_06772_),
    .A2_N(_06773_),
    .B1(_06760_),
    .B2(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__a21oi_2 _12425_ (.A1(_06748_),
    .A2(_06360_),
    .B1(_06362_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_2 _12426_ (.A(_06398_),
    .B(_06751_),
    .Y(_06779_));
 sky130_fd_sc_hd__or2b_1 _12427_ (.A(_06390_),
    .B_N(_06756_),
    .X(_06780_));
 sky130_fd_sc_hd__clkbuf_4 _12428_ (.A(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__a41o_1 _12429_ (.A1(_06363_),
    .A2(_06753_),
    .A3(_06781_),
    .A4(_06766_),
    .B1(_06358_),
    .X(_06782_));
 sky130_fd_sc_hd__a21oi_1 _12430_ (.A1(_06778_),
    .A2(_06779_),
    .B1(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__nand2b_4 _12431_ (.A_N(_06379_),
    .B(_06756_),
    .Y(_06784_));
 sky130_fd_sc_hd__a21oi_1 _12432_ (.A1(_06748_),
    .A2(_06784_),
    .B1(_06363_),
    .Y(_06785_));
 sky130_fd_sc_hd__nand3b_4 _12433_ (.A_N(_06756_),
    .B(_06379_),
    .C(_06390_),
    .Y(_06786_));
 sky130_fd_sc_hd__a31o_1 _12434_ (.A1(_06363_),
    .A2(_06781_),
    .A3(_06786_),
    .B1(_06401_),
    .X(_06787_));
 sky130_fd_sc_hd__o21ai_1 _12435_ (.A1(_06785_),
    .A2(_06787_),
    .B1(\sinegen0.read_ptr[6] ),
    .Y(_06788_));
 sky130_fd_sc_hd__o221a_1 _12436_ (.A1(_06747_),
    .A2(_06777_),
    .B1(_06783_),
    .B2(_06788_),
    .C1(_06405_),
    .X(_06789_));
 sky130_fd_sc_hd__a211oi_2 _12437_ (.A1(_06370_),
    .A2(_06771_),
    .B1(_06789_),
    .C1(_06357_),
    .Y(_06790_));
 sky130_fd_sc_hd__a21oi_1 _12438_ (.A1(_06611_),
    .A2(_06746_),
    .B1(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__buf_8 _12439_ (.A(_06643_),
    .X(_06792_));
 sky130_fd_sc_hd__buf_12 _12440_ (.A(_06621_),
    .X(_06793_));
 sky130_fd_sc_hd__mux4_2 _12441_ (.A0(\fifo0.fifo_store[96][13] ),
    .A1(\fifo0.fifo_store[97][13] ),
    .A2(\fifo0.fifo_store[98][13] ),
    .A3(\fifo0.fifo_store[99][13] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_06794_));
 sky130_fd_sc_hd__buf_12 _12442_ (.A(_06450_),
    .X(_06795_));
 sky130_fd_sc_hd__mux4_1 _12443_ (.A0(\fifo0.fifo_store[100][13] ),
    .A1(\fifo0.fifo_store[101][13] ),
    .A2(\fifo0.fifo_store[102][13] ),
    .A3(\fifo0.fifo_store[103][13] ),
    .S0(_06795_),
    .S1(_06504_),
    .X(_06796_));
 sky130_fd_sc_hd__buf_12 _12444_ (.A(_06440_),
    .X(_06797_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(_06794_),
    .A1(_06796_),
    .S(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__mux4_1 _12446_ (.A0(\fifo0.fifo_store[104][13] ),
    .A1(\fifo0.fifo_store[105][13] ),
    .A2(\fifo0.fifo_store[106][13] ),
    .A3(\fifo0.fifo_store[107][13] ),
    .S0(_06693_),
    .S1(_06579_),
    .X(_06799_));
 sky130_fd_sc_hd__or2_1 _12447_ (.A(_06624_),
    .B(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__buf_8 _12448_ (.A(_06673_),
    .X(_06801_));
 sky130_fd_sc_hd__mux4_1 _12449_ (.A0(\fifo0.fifo_store[108][13] ),
    .A1(\fifo0.fifo_store[109][13] ),
    .A2(\fifo0.fifo_store[110][13] ),
    .A3(\fifo0.fifo_store[111][13] ),
    .S0(_06801_),
    .S1(_06421_),
    .X(_06802_));
 sky130_fd_sc_hd__o21a_1 _12450_ (.A1(_06681_),
    .A2(_06802_),
    .B1(_06630_),
    .X(_06803_));
 sky130_fd_sc_hd__buf_12 _12451_ (.A(_06641_),
    .X(_06804_));
 sky130_fd_sc_hd__a221o_1 _12452_ (.A1(_06793_),
    .A2(_06798_),
    .B1(_06800_),
    .B2(_06803_),
    .C1(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__or2_1 _12453_ (.A(_06612_),
    .B(\fifo0.fifo_store[119][13] ),
    .X(_06806_));
 sky130_fd_sc_hd__o21a_1 _12454_ (.A1(_06435_),
    .A2(\fifo0.fifo_store[118][13] ),
    .B1(_06615_),
    .X(_06807_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\fifo0.fifo_store[116][13] ),
    .A1(\fifo0.fifo_store[117][13] ),
    .S(_06689_),
    .X(_06808_));
 sky130_fd_sc_hd__a221o_1 _12456_ (.A1(_06806_),
    .A2(_06807_),
    .B1(_06808_),
    .B2(_06425_),
    .C1(_06477_),
    .X(_06809_));
 sky130_fd_sc_hd__clkbuf_16 _12457_ (.A(_06520_),
    .X(_06810_));
 sky130_fd_sc_hd__buf_12 _12458_ (.A(_06627_),
    .X(_06811_));
 sky130_fd_sc_hd__mux4_1 _12459_ (.A0(\fifo0.fifo_store[112][13] ),
    .A1(\fifo0.fifo_store[113][13] ),
    .A2(\fifo0.fifo_store[114][13] ),
    .A3(\fifo0.fifo_store[115][13] ),
    .S0(_06810_),
    .S1(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__or2_1 _12460_ (.A(_06599_),
    .B(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_16 _12461_ (.A(_06634_),
    .X(_06814_));
 sky130_fd_sc_hd__mux4_1 _12462_ (.A0(\fifo0.fifo_store[124][13] ),
    .A1(\fifo0.fifo_store[125][13] ),
    .A2(\fifo0.fifo_store[126][13] ),
    .A3(\fifo0.fifo_store[127][13] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_06815_));
 sky130_fd_sc_hd__mux4_2 _12463_ (.A0(\fifo0.fifo_store[120][13] ),
    .A1(\fifo0.fifo_store[121][13] ),
    .A2(\fifo0.fifo_store[122][13] ),
    .A3(\fifo0.fifo_store[123][13] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_06816_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(_06623_),
    .B(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__o211a_1 _12465_ (.A1(_06814_),
    .A2(_06815_),
    .B1(_06817_),
    .C1(_06664_),
    .X(_06818_));
 sky130_fd_sc_hd__a311o_1 _12466_ (.A1(_06793_),
    .A2(_06809_),
    .A3(_06813_),
    .B1(_06494_),
    .C1(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__mux4_1 _12467_ (.A0(\fifo0.fifo_store[76][13] ),
    .A1(\fifo0.fifo_store[77][13] ),
    .A2(\fifo0.fifo_store[78][13] ),
    .A3(\fifo0.fifo_store[79][13] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_06820_));
 sky130_fd_sc_hd__mux4_1 _12468_ (.A0(\fifo0.fifo_store[72][13] ),
    .A1(\fifo0.fifo_store[73][13] ),
    .A2(\fifo0.fifo_store[74][13] ),
    .A3(\fifo0.fifo_store[75][13] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_06821_));
 sky130_fd_sc_hd__or2_1 _12469_ (.A(_06623_),
    .B(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__o211a_2 _12470_ (.A1(_06814_),
    .A2(_06820_),
    .B1(_06822_),
    .C1(_06630_),
    .X(_06823_));
 sky130_fd_sc_hd__buf_8 _12471_ (.A(_06683_),
    .X(_06824_));
 sky130_fd_sc_hd__mux4_1 _12472_ (.A0(\fifo0.fifo_store[64][13] ),
    .A1(\fifo0.fifo_store[65][13] ),
    .A2(\fifo0.fifo_store[66][13] ),
    .A3(\fifo0.fifo_store[67][13] ),
    .S0(_06549_),
    .S1(_06615_),
    .X(_06825_));
 sky130_fd_sc_hd__or2b_1 _12473_ (.A(\fifo0.fifo_store[71][13] ),
    .B_N(_06521_),
    .X(_06826_));
 sky130_fd_sc_hd__o21a_1 _12474_ (.A1(_06536_),
    .A2(\fifo0.fifo_store[70][13] ),
    .B1(_06690_),
    .X(_06827_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(\fifo0.fifo_store[68][13] ),
    .A1(\fifo0.fifo_store[69][13] ),
    .S(_06544_),
    .X(_06828_));
 sky130_fd_sc_hd__buf_8 _12476_ (.A(_06424_),
    .X(_06829_));
 sky130_fd_sc_hd__a221o_1 _12477_ (.A1(_06826_),
    .A2(_06827_),
    .B1(_06828_),
    .B2(_06829_),
    .C1(_06634_),
    .X(_06830_));
 sky130_fd_sc_hd__o211a_1 _12478_ (.A1(_06824_),
    .A2(_06825_),
    .B1(_06830_),
    .C1(_06735_),
    .X(_06831_));
 sky130_fd_sc_hd__mux4_1 _12479_ (.A0(\fifo0.fifo_store[80][13] ),
    .A1(\fifo0.fifo_store[81][13] ),
    .A2(\fifo0.fifo_store[82][13] ),
    .A3(\fifo0.fifo_store[83][13] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_06832_));
 sky130_fd_sc_hd__mux4_1 _12480_ (.A0(\fifo0.fifo_store[84][13] ),
    .A1(\fifo0.fifo_store[85][13] ),
    .A2(\fifo0.fifo_store[86][13] ),
    .A3(\fifo0.fifo_store[87][13] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_06833_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(_06832_),
    .A1(_06833_),
    .S(_06447_),
    .X(_06834_));
 sky130_fd_sc_hd__mux4_1 _12482_ (.A0(\fifo0.fifo_store[88][13] ),
    .A1(\fifo0.fifo_store[89][13] ),
    .A2(\fifo0.fifo_store[90][13] ),
    .A3(\fifo0.fifo_store[91][13] ),
    .S0(_06673_),
    .S1(_06420_),
    .X(_06835_));
 sky130_fd_sc_hd__or2_1 _12483_ (.A(_06683_),
    .B(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__mux4_2 _12484_ (.A0(\fifo0.fifo_store[92][13] ),
    .A1(\fifo0.fifo_store[93][13] ),
    .A2(\fifo0.fifo_store[94][13] ),
    .A3(\fifo0.fifo_store[95][13] ),
    .S0(_06717_),
    .S1(_06718_),
    .X(_06837_));
 sky130_fd_sc_hd__o21a_1 _12485_ (.A1(_06680_),
    .A2(_06837_),
    .B1(_06663_),
    .X(_06838_));
 sky130_fd_sc_hd__a221o_1 _12486_ (.A1(_06735_),
    .A2(_06834_),
    .B1(_06836_),
    .B2(_06838_),
    .C1(_06743_),
    .X(_06839_));
 sky130_fd_sc_hd__o311a_1 _12487_ (.A1(_06804_),
    .A2(_06823_),
    .A3(_06831_),
    .B1(_06839_),
    .C1(_06677_),
    .X(_06840_));
 sky130_fd_sc_hd__a311o_4 _12488_ (.A1(_06792_),
    .A2(_06805_),
    .A3(_06819_),
    .B1(_06604_),
    .C1(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__or2_1 _12489_ (.A(_06527_),
    .B(\fifo0.fifo_store[4][13] ),
    .X(_06842_));
 sky130_fd_sc_hd__o211a_1 _12490_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[5][13] ),
    .B1(_06842_),
    .C1(_06650_),
    .X(_06843_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\fifo0.fifo_store[6][13] ),
    .A1(\fifo0.fifo_store[7][13] ),
    .S(_06617_),
    .X(_06844_));
 sky130_fd_sc_hd__a21o_1 _12492_ (.A1(_06648_),
    .A2(_06844_),
    .B1(_06476_),
    .X(_06845_));
 sky130_fd_sc_hd__mux4_1 _12493_ (.A0(\fifo0.fifo_store[0][13] ),
    .A1(\fifo0.fifo_store[1][13] ),
    .A2(\fifo0.fifo_store[2][13] ),
    .A3(\fifo0.fifo_store[3][13] ),
    .S0(_06479_),
    .S1(_06811_),
    .X(_06846_));
 sky130_fd_sc_hd__o221a_1 _12494_ (.A1(_06843_),
    .A2(_06845_),
    .B1(_06846_),
    .B2(_06599_),
    .C1(_06621_),
    .X(_06847_));
 sky130_fd_sc_hd__buf_8 _12495_ (.A(_06657_),
    .X(_06848_));
 sky130_fd_sc_hd__mux4_2 _12496_ (.A0(\fifo0.fifo_store[8][13] ),
    .A1(\fifo0.fifo_store[9][13] ),
    .A2(\fifo0.fifo_store[10][13] ),
    .A3(\fifo0.fifo_store[11][13] ),
    .S0(_06848_),
    .S1(_06511_),
    .X(_06849_));
 sky130_fd_sc_hd__mux4_2 _12497_ (.A0(\fifo0.fifo_store[12][13] ),
    .A1(\fifo0.fifo_store[13][13] ),
    .A2(\fifo0.fifo_store[14][13] ),
    .A3(\fifo0.fifo_store[15][13] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_06850_));
 sky130_fd_sc_hd__or2_1 _12498_ (.A(_06660_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__o211a_1 _12499_ (.A1(_06656_),
    .A2(_06849_),
    .B1(_06851_),
    .C1(_06630_),
    .X(_06852_));
 sky130_fd_sc_hd__mux4_1 _12500_ (.A0(\fifo0.fifo_store[24][13] ),
    .A1(\fifo0.fifo_store[25][13] ),
    .A2(\fifo0.fifo_store[26][13] ),
    .A3(\fifo0.fifo_store[27][13] ),
    .S0(_06657_),
    .S1(_06578_),
    .X(_06853_));
 sky130_fd_sc_hd__or2_1 _12501_ (.A(_06623_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__mux4_1 _12502_ (.A0(\fifo0.fifo_store[28][13] ),
    .A1(\fifo0.fifo_store[29][13] ),
    .A2(\fifo0.fifo_store[30][13] ),
    .A3(\fifo0.fifo_store[31][13] ),
    .S0(_06673_),
    .S1(_06614_),
    .X(_06855_));
 sky130_fd_sc_hd__o21a_1 _12503_ (.A1(_06680_),
    .A2(_06855_),
    .B1(_06461_),
    .X(_06856_));
 sky130_fd_sc_hd__mux4_1 _12504_ (.A0(\fifo0.fifo_store[16][13] ),
    .A1(\fifo0.fifo_store[17][13] ),
    .A2(\fifo0.fifo_store[18][13] ),
    .A3(\fifo0.fifo_store[19][13] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_06857_));
 sky130_fd_sc_hd__or2_1 _12505_ (.A(_06655_),
    .B(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__mux4_1 _12506_ (.A0(\fifo0.fifo_store[20][13] ),
    .A1(\fifo0.fifo_store[21][13] ),
    .A2(\fifo0.fifo_store[22][13] ),
    .A3(\fifo0.fifo_store[23][13] ),
    .S0(_06548_),
    .S1(_06703_),
    .X(_06859_));
 sky130_fd_sc_hd__o21a_1 _12507_ (.A1(_06680_),
    .A2(_06859_),
    .B1(_06466_),
    .X(_06860_));
 sky130_fd_sc_hd__a221o_1 _12508_ (.A1(_06854_),
    .A2(_06856_),
    .B1(_06858_),
    .B2(_06860_),
    .C1(_06743_),
    .X(_06861_));
 sky130_fd_sc_hd__o311a_4 _12509_ (.A1(_06589_),
    .A2(_06847_),
    .A3(_06852_),
    .B1(_06677_),
    .C1(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__or2_1 _12510_ (.A(_06434_),
    .B(\fifo0.fifo_store[52][13] ),
    .X(_06863_));
 sky130_fd_sc_hd__o211a_1 _12511_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[53][13] ),
    .B1(_06863_),
    .C1(_06728_),
    .X(_06864_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(\fifo0.fifo_store[54][13] ),
    .A1(\fifo0.fifo_store[55][13] ),
    .S(_06710_),
    .X(_06865_));
 sky130_fd_sc_hd__a21o_1 _12513_ (.A1(_06691_),
    .A2(_06865_),
    .B1(_06660_),
    .X(_06866_));
 sky130_fd_sc_hd__mux4_1 _12514_ (.A0(\fifo0.fifo_store[48][13] ),
    .A1(\fifo0.fifo_store[49][13] ),
    .A2(\fifo0.fifo_store[50][13] ),
    .A3(\fifo0.fifo_store[51][13] ),
    .S0(_06487_),
    .S1(_06489_),
    .X(_06867_));
 sky130_fd_sc_hd__clkbuf_16 _12515_ (.A(_06466_),
    .X(_06868_));
 sky130_fd_sc_hd__o221a_1 _12516_ (.A1(_06864_),
    .A2(_06866_),
    .B1(_06867_),
    .B2(_06624_),
    .C1(_06868_),
    .X(_06869_));
 sky130_fd_sc_hd__buf_8 _12517_ (.A(_06548_),
    .X(_06870_));
 sky130_fd_sc_hd__mux4_1 _12518_ (.A0(\fifo0.fifo_store[56][13] ),
    .A1(\fifo0.fifo_store[57][13] ),
    .A2(\fifo0.fifo_store[58][13] ),
    .A3(\fifo0.fifo_store[59][13] ),
    .S0(_06870_),
    .S1(_06615_),
    .X(_06871_));
 sky130_fd_sc_hd__mux4_1 _12519_ (.A0(\fifo0.fifo_store[60][13] ),
    .A1(\fifo0.fifo_store[61][13] ),
    .A2(\fifo0.fifo_store[62][13] ),
    .A3(\fifo0.fifo_store[63][13] ),
    .S0(_06657_),
    .S1(_06578_),
    .X(_06872_));
 sky130_fd_sc_hd__or2_1 _12520_ (.A(_06634_),
    .B(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__o211a_1 _12521_ (.A1(_06824_),
    .A2(_06871_),
    .B1(_06873_),
    .C1(_06664_),
    .X(_06874_));
 sky130_fd_sc_hd__mux4_1 _12522_ (.A0(\fifo0.fifo_store[40][13] ),
    .A1(\fifo0.fifo_store[41][13] ),
    .A2(\fifo0.fifo_store[42][13] ),
    .A3(\fifo0.fifo_store[43][13] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_06875_));
 sky130_fd_sc_hd__or2_1 _12523_ (.A(_06655_),
    .B(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__mux4_1 _12524_ (.A0(\fifo0.fifo_store[44][13] ),
    .A1(\fifo0.fifo_store[45][13] ),
    .A2(\fifo0.fifo_store[46][13] ),
    .A3(\fifo0.fifo_store[47][13] ),
    .S0(_06548_),
    .S1(_06614_),
    .X(_06877_));
 sky130_fd_sc_hd__o21a_1 _12525_ (.A1(_06680_),
    .A2(_06877_),
    .B1(_06663_),
    .X(_06878_));
 sky130_fd_sc_hd__mux4_1 _12526_ (.A0(\fifo0.fifo_store[32][13] ),
    .A1(\fifo0.fifo_store[33][13] ),
    .A2(\fifo0.fifo_store[34][13] ),
    .A3(\fifo0.fifo_store[35][13] ),
    .S0(_06673_),
    .S1(_06420_),
    .X(_06879_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(_06655_),
    .B(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__mux4_1 _12528_ (.A0(\fifo0.fifo_store[36][13] ),
    .A1(\fifo0.fifo_store[37][13] ),
    .A2(\fifo0.fifo_store[38][13] ),
    .A3(\fifo0.fifo_store[39][13] ),
    .S0(_06717_),
    .S1(_06703_),
    .X(_06881_));
 sky130_fd_sc_hd__o21a_1 _12529_ (.A1(_06680_),
    .A2(_06881_),
    .B1(_06466_),
    .X(_06882_));
 sky130_fd_sc_hd__a221o_1 _12530_ (.A1(_06876_),
    .A2(_06878_),
    .B1(_06880_),
    .B2(_06882_),
    .C1(_06641_),
    .X(_06883_));
 sky130_fd_sc_hd__o311a_4 _12531_ (.A1(_06679_),
    .A2(_06869_),
    .A3(_06874_),
    .B1(_06883_),
    .C1(_06643_),
    .X(_06884_));
 sky130_fd_sc_hd__o31a_1 _12532_ (.A1(_00006_),
    .A2(_06862_),
    .A3(_06884_),
    .B1(_06357_),
    .X(_06885_));
 sky130_fd_sc_hd__a21oi_2 _12533_ (.A1(_06364_),
    .A2(_06365_),
    .B1(_06366_),
    .Y(_06886_));
 sky130_fd_sc_hd__a21o_1 _12534_ (.A1(_06391_),
    .A2(_06360_),
    .B1(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__nor2_1 _12535_ (.A(_06361_),
    .B(_06775_),
    .Y(_06888_));
 sky130_fd_sc_hd__a21oi_1 _12536_ (.A1(_06396_),
    .A2(_06887_),
    .B1(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__nor2_1 _12537_ (.A(_06391_),
    .B(_06380_),
    .Y(_06890_));
 sky130_fd_sc_hd__a21oi_4 _12538_ (.A1(_06390_),
    .A2(_06379_),
    .B1(_06376_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_1 _12539_ (.A(_06366_),
    .B(_06365_),
    .Y(_06892_));
 sky130_fd_sc_hd__a21o_1 _12540_ (.A1(_06892_),
    .A2(_06386_),
    .B1(_06362_),
    .X(_06893_));
 sky130_fd_sc_hd__o31a_1 _12541_ (.A1(_06382_),
    .A2(_06890_),
    .A3(_06891_),
    .B1(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__a21oi_1 _12542_ (.A1(_06397_),
    .A2(_06781_),
    .B1(_06751_),
    .Y(_06895_));
 sky130_fd_sc_hd__nor2_1 _12543_ (.A(_06888_),
    .B(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__nand2_1 _12544_ (.A(_06379_),
    .B(_06756_),
    .Y(_06897_));
 sky130_fd_sc_hd__or2_1 _12545_ (.A(_06395_),
    .B(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__and3_2 _12546_ (.A(_06384_),
    .B(_06753_),
    .C(_06765_),
    .X(_06899_));
 sky130_fd_sc_hd__o2bb2a_1 _12547_ (.A1_N(_06898_),
    .A2_N(_06899_),
    .B1(_06897_),
    .B2(_06775_),
    .X(_06900_));
 sky130_fd_sc_hd__mux4_1 _12548_ (.A0(_06889_),
    .A1(_06894_),
    .A2(_06896_),
    .A3(_06900_),
    .S0(_06404_),
    .S1(_06402_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_4 _12549_ (.A(_06373_),
    .X(_06902_));
 sky130_fd_sc_hd__a21oi_1 _12550_ (.A1(_06748_),
    .A2(_06751_),
    .B1(_06396_),
    .Y(_06903_));
 sky130_fd_sc_hd__a21oi_1 _12551_ (.A1(_06386_),
    .A2(_06786_),
    .B1(_06378_),
    .Y(_06904_));
 sky130_fd_sc_hd__or3b_1 _12552_ (.A(_06364_),
    .B(_06365_),
    .C_N(_06366_),
    .X(_06905_));
 sky130_fd_sc_hd__a32o_1 _12553_ (.A1(_06397_),
    .A2(_06384_),
    .A3(_06905_),
    .B1(_06784_),
    .B2(_06891_),
    .X(_06906_));
 sky130_fd_sc_hd__nand2_1 _12554_ (.A(_06902_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__o311a_1 _12555_ (.A1(_06902_),
    .A2(_06903_),
    .A3(_06904_),
    .B1(_06907_),
    .C1(_06404_),
    .X(_06908_));
 sky130_fd_sc_hd__a211oi_1 _12556_ (.A1(_06363_),
    .A2(_06887_),
    .B1(_06760_),
    .C1(_06762_),
    .Y(_06909_));
 sky130_fd_sc_hd__and2b_2 _12557_ (.A_N(\sinegen0.read_ptr[5] ),
    .B(\sinegen0.read_ptr[4] ),
    .X(_06910_));
 sky130_fd_sc_hd__and2b_1 _12558_ (.A_N(_06376_),
    .B(_06379_),
    .X(_06911_));
 sky130_fd_sc_hd__o21bai_4 _12559_ (.A1(_06366_),
    .A2(_06365_),
    .B1_N(_06376_),
    .Y(_06912_));
 sky130_fd_sc_hd__a21oi_1 _12560_ (.A1(_06391_),
    .A2(_06750_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__a211o_1 _12561_ (.A1(_06766_),
    .A2(_06911_),
    .B1(_06888_),
    .C1(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__a221o_1 _12562_ (.A1(_06369_),
    .A2(_06909_),
    .B1(_06910_),
    .B2(_06914_),
    .C1(\sinegen0.read_ptr[6] ),
    .X(_06915_));
 sky130_fd_sc_hd__o221a_1 _12563_ (.A1(_06769_),
    .A2(_06901_),
    .B1(_06908_),
    .B2(_06915_),
    .C1(net23),
    .X(_06916_));
 sky130_fd_sc_hd__a21oi_1 _12564_ (.A1(_06841_),
    .A2(_06885_),
    .B1(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__buf_4 _12565_ (.A(net23),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_4 _12566_ (.A(\sinegen0.read_ptr[6] ),
    .X(_06919_));
 sky130_fd_sc_hd__nor2_1 _12567_ (.A(_06748_),
    .B(_06751_),
    .Y(_06920_));
 sky130_fd_sc_hd__a32o_1 _12568_ (.A1(_06397_),
    .A2(_06361_),
    .A3(_06781_),
    .B1(_06383_),
    .B2(_06388_),
    .X(_06921_));
 sky130_fd_sc_hd__nor2_4 _12569_ (.A(_06376_),
    .B(_06364_),
    .Y(_06922_));
 sky130_fd_sc_hd__xnor2_4 _12570_ (.A(_06390_),
    .B(_06756_),
    .Y(_06923_));
 sky130_fd_sc_hd__or2_1 _12571_ (.A(_06390_),
    .B(_06756_),
    .X(_06924_));
 sky130_fd_sc_hd__and3_1 _12572_ (.A(_06362_),
    .B(_06924_),
    .C(_06784_),
    .X(_06925_));
 sky130_fd_sc_hd__a21o_1 _12573_ (.A1(_06922_),
    .A2(_06923_),
    .B1(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__or2_1 _12574_ (.A(_06376_),
    .B(_06365_),
    .X(_06927_));
 sky130_fd_sc_hd__and2_1 _12575_ (.A(_06753_),
    .B(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__mux4_1 _12576_ (.A0(_06920_),
    .A1(_06921_),
    .A2(_06926_),
    .A3(_06928_),
    .S0(_06369_),
    .S1(_06402_),
    .X(_06929_));
 sky130_fd_sc_hd__and3_1 _12577_ (.A(_06395_),
    .B(_06361_),
    .C(_06781_),
    .X(_06930_));
 sky130_fd_sc_hd__o21ai_1 _12578_ (.A1(_06925_),
    .A2(_06930_),
    .B1(_06902_),
    .Y(_06931_));
 sky130_fd_sc_hd__o211a_1 _12579_ (.A1(_06778_),
    .A2(_06782_),
    .B1(_06931_),
    .C1(_06404_),
    .X(_06932_));
 sky130_fd_sc_hd__a21o_1 _12580_ (.A1(_06361_),
    .A2(_06781_),
    .B1(_06395_),
    .X(_06933_));
 sky130_fd_sc_hd__nand2_1 _12581_ (.A(_06911_),
    .B(_06923_),
    .Y(_06934_));
 sky130_fd_sc_hd__o311a_1 _12582_ (.A1(_06377_),
    .A2(_06890_),
    .A3(_06759_),
    .B1(_06372_),
    .C1(_06401_),
    .X(_06935_));
 sky130_fd_sc_hd__a311o_1 _12583_ (.A1(_06902_),
    .A2(_06933_),
    .A3(_06934_),
    .B1(_06935_),
    .C1(_06404_),
    .X(_06936_));
 sky130_fd_sc_hd__nand2_1 _12584_ (.A(_06747_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__o22a_1 _12585_ (.A1(_06919_),
    .A2(_06929_),
    .B1(_06932_),
    .B2(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_16 _12586_ (.A(_06701_),
    .X(_06939_));
 sky130_fd_sc_hd__mux4_2 _12587_ (.A0(\fifo0.fifo_store[96][12] ),
    .A1(\fifo0.fifo_store[97][12] ),
    .A2(\fifo0.fifo_store[98][12] ),
    .A3(\fifo0.fifo_store[99][12] ),
    .S0(_06693_),
    .S1(_06579_),
    .X(_06940_));
 sky130_fd_sc_hd__mux4_1 _12588_ (.A0(\fifo0.fifo_store[100][12] ),
    .A1(\fifo0.fifo_store[101][12] ),
    .A2(\fifo0.fifo_store[102][12] ),
    .A3(\fifo0.fifo_store[103][12] ),
    .S0(_06625_),
    .S1(_06579_),
    .X(_06941_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(_06940_),
    .A1(_06941_),
    .S(_06448_),
    .X(_06942_));
 sky130_fd_sc_hd__mux4_1 _12590_ (.A0(\fifo0.fifo_store[104][12] ),
    .A1(\fifo0.fifo_store[105][12] ),
    .A2(\fifo0.fifo_store[106][12] ),
    .A3(\fifo0.fifo_store[107][12] ),
    .S0(_06514_),
    .S1(_06615_),
    .X(_06943_));
 sky130_fd_sc_hd__or2_1 _12591_ (.A(_06824_),
    .B(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__buf_8 _12592_ (.A(_06721_),
    .X(_06945_));
 sky130_fd_sc_hd__buf_12 _12593_ (.A(_06513_),
    .X(_06946_));
 sky130_fd_sc_hd__mux4_1 _12594_ (.A0(\fifo0.fifo_store[108][12] ),
    .A1(\fifo0.fifo_store[109][12] ),
    .A2(\fifo0.fifo_store[110][12] ),
    .A3(\fifo0.fifo_store[111][12] ),
    .S0(_06946_),
    .S1(_06648_),
    .X(_06947_));
 sky130_fd_sc_hd__o21a_1 _12595_ (.A1(_06945_),
    .A2(_06947_),
    .B1(_06664_),
    .X(_06948_));
 sky130_fd_sc_hd__a221o_1 _12596_ (.A1(_06939_),
    .A2(_06942_),
    .B1(_06944_),
    .B2(_06948_),
    .C1(_06804_),
    .X(_06949_));
 sky130_fd_sc_hd__or2_1 _12597_ (.A(_06612_),
    .B(\fifo0.fifo_store[119][12] ),
    .X(_06950_));
 sky130_fd_sc_hd__buf_12 _12598_ (.A(_06600_),
    .X(_06951_));
 sky130_fd_sc_hd__o21a_1 _12599_ (.A1(_06951_),
    .A2(\fifo0.fifo_store[118][12] ),
    .B1(_06691_),
    .X(_06952_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(\fifo0.fifo_store[116][12] ),
    .A1(\fifo0.fifo_store[117][12] ),
    .S(_06576_),
    .X(_06953_));
 sky130_fd_sc_hd__buf_8 _12601_ (.A(_06424_),
    .X(_06954_));
 sky130_fd_sc_hd__a221o_1 _12602_ (.A1(_06950_),
    .A2(_06952_),
    .B1(_06953_),
    .B2(_06954_),
    .C1(_06681_),
    .X(_06955_));
 sky130_fd_sc_hd__buf_8 _12603_ (.A(_06673_),
    .X(_06956_));
 sky130_fd_sc_hd__mux4_1 _12604_ (.A0(\fifo0.fifo_store[112][12] ),
    .A1(\fifo0.fifo_store[113][12] ),
    .A2(\fifo0.fifo_store[114][12] ),
    .A3(\fifo0.fifo_store[115][12] ),
    .S0(_06956_),
    .S1(_06421_),
    .X(_06957_));
 sky130_fd_sc_hd__or2_1 _12605_ (.A(_06656_),
    .B(_06957_),
    .X(_06958_));
 sky130_fd_sc_hd__buf_12 _12606_ (.A(_06513_),
    .X(_06959_));
 sky130_fd_sc_hd__mux4_1 _12607_ (.A0(\fifo0.fifo_store[124][12] ),
    .A1(\fifo0.fifo_store[125][12] ),
    .A2(\fifo0.fifo_store[126][12] ),
    .A3(\fifo0.fifo_store[127][12] ),
    .S0(_06959_),
    .S1(_06648_),
    .X(_06960_));
 sky130_fd_sc_hd__mux4_1 _12608_ (.A0(\fifo0.fifo_store[120][12] ),
    .A1(\fifo0.fifo_store[121][12] ),
    .A2(\fifo0.fifo_store[122][12] ),
    .A3(\fifo0.fifo_store[123][12] ),
    .S0(_06717_),
    .S1(_06718_),
    .X(_06961_));
 sky130_fd_sc_hd__or2_1 _12609_ (.A(_06683_),
    .B(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__o211a_1 _12610_ (.A1(_06681_),
    .A2(_06960_),
    .B1(_06962_),
    .C1(_06686_),
    .X(_06963_));
 sky130_fd_sc_hd__a311o_1 _12611_ (.A1(_06939_),
    .A2(_06955_),
    .A3(_06958_),
    .B1(_06679_),
    .C1(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__buf_12 _12612_ (.A(_06604_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_16 _12613_ (.A(_06641_),
    .X(_06966_));
 sky130_fd_sc_hd__mux4_1 _12614_ (.A0(\fifo0.fifo_store[76][12] ),
    .A1(\fifo0.fifo_store[77][12] ),
    .A2(\fifo0.fifo_store[78][12] ),
    .A3(\fifo0.fifo_store[79][12] ),
    .S0(_06946_),
    .S1(_06691_),
    .X(_06967_));
 sky130_fd_sc_hd__mux4_1 _12615_ (.A0(\fifo0.fifo_store[72][12] ),
    .A1(\fifo0.fifo_store[73][12] ),
    .A2(\fifo0.fifo_store[74][12] ),
    .A3(\fifo0.fifo_store[75][12] ),
    .S0(_06513_),
    .S1(_06647_),
    .X(_06968_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(_06730_),
    .B(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__o211a_1 _12617_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_06969_),
    .C1(_06686_),
    .X(_06970_));
 sky130_fd_sc_hd__buf_12 _12618_ (.A(_06711_),
    .X(_06971_));
 sky130_fd_sc_hd__mux4_2 _12619_ (.A0(\fifo0.fifo_store[64][12] ),
    .A1(\fifo0.fifo_store[65][12] ),
    .A2(\fifo0.fifo_store[66][12] ),
    .A3(\fifo0.fifo_store[67][12] ),
    .S0(_06416_),
    .S1(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_12 _12620_ (.A(_06673_),
    .X(_06973_));
 sky130_fd_sc_hd__or2b_1 _12621_ (.A(\fifo0.fifo_store[71][12] ),
    .B_N(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__clkbuf_16 _12622_ (.A(_06470_),
    .X(_06975_));
 sky130_fd_sc_hd__o21a_1 _12623_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[70][12] ),
    .B1(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__buf_12 _12624_ (.A(_06433_),
    .X(_06977_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(\fifo0.fifo_store[68][12] ),
    .A1(\fifo0.fifo_store[69][12] ),
    .S(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__a221o_1 _12626_ (.A1(_06974_),
    .A2(_06976_),
    .B1(_06978_),
    .B2(_06699_),
    .C1(_06721_),
    .X(_06979_));
 sky130_fd_sc_hd__o211a_1 _12627_ (.A1(_06688_),
    .A2(_06972_),
    .B1(_06979_),
    .C1(_06701_),
    .X(_06980_));
 sky130_fd_sc_hd__mux4_1 _12628_ (.A0(\fifo0.fifo_store[80][12] ),
    .A1(\fifo0.fifo_store[81][12] ),
    .A2(\fifo0.fifo_store[82][12] ),
    .A3(\fifo0.fifo_store[83][12] ),
    .S0(_06717_),
    .S1(_06703_),
    .X(_06981_));
 sky130_fd_sc_hd__mux4_1 _12629_ (.A0(\fifo0.fifo_store[84][12] ),
    .A1(\fifo0.fifo_store[85][12] ),
    .A2(\fifo0.fifo_store[86][12] ),
    .A3(\fifo0.fifo_store[87][12] ),
    .S0(_06717_),
    .S1(_06703_),
    .X(_06982_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(_06981_),
    .A1(_06982_),
    .S(_06484_),
    .X(_06983_));
 sky130_fd_sc_hd__buf_12 _12631_ (.A(_06419_),
    .X(_06984_));
 sky130_fd_sc_hd__mux4_1 _12632_ (.A0(\fifo0.fifo_store[88][12] ),
    .A1(\fifo0.fifo_store[89][12] ),
    .A2(\fifo0.fifo_store[90][12] ),
    .A3(\fifo0.fifo_store[91][12] ),
    .S0(_06415_),
    .S1(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__or2_1 _12633_ (.A(_06531_),
    .B(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__mux4_2 _12634_ (.A0(\fifo0.fifo_store[92][12] ),
    .A1(\fifo0.fifo_store[93][12] ),
    .A2(\fifo0.fifo_store[94][12] ),
    .A3(\fifo0.fifo_store[95][12] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_06987_));
 sky130_fd_sc_hd__o21a_1 _12635_ (.A1(_06709_),
    .A2(_06987_),
    .B1(_06713_),
    .X(_06988_));
 sky130_fd_sc_hd__a221o_1 _12636_ (.A1(_06701_),
    .A2(_06983_),
    .B1(_06986_),
    .B2(_06988_),
    .C1(_06743_),
    .X(_06989_));
 sky130_fd_sc_hd__o311a_1 _12637_ (.A1(_06966_),
    .A2(_06970_),
    .A3(_06980_),
    .B1(_06989_),
    .C1(_06498_),
    .X(_06990_));
 sky130_fd_sc_hd__a311oi_4 _12638_ (.A1(_06792_),
    .A2(_06949_),
    .A3(_06964_),
    .B1(_06965_),
    .C1(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__buf_12 _12639_ (.A(_00006_),
    .X(_06992_));
 sky130_fd_sc_hd__buf_6 _12640_ (.A(_06412_),
    .X(_06993_));
 sky130_fd_sc_hd__or2_1 _12641_ (.A(_06479_),
    .B(\fifo0.fifo_store[4][12] ),
    .X(_06994_));
 sky130_fd_sc_hd__o211a_1 _12642_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[5][12] ),
    .B1(_06994_),
    .C1(_06699_),
    .X(_06995_));
 sky130_fd_sc_hd__buf_12 _12643_ (.A(_06528_),
    .X(_06996_));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(\fifo0.fifo_store[6][12] ),
    .A1(\fifo0.fifo_store[7][12] ),
    .S(_06697_),
    .X(_06997_));
 sky130_fd_sc_hd__a21o_1 _12645_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_06680_),
    .X(_06998_));
 sky130_fd_sc_hd__mux4_1 _12646_ (.A0(\fifo0.fifo_store[0][12] ),
    .A1(\fifo0.fifo_store[1][12] ),
    .A2(\fifo0.fifo_store[2][12] ),
    .A3(\fifo0.fifo_store[3][12] ),
    .S0(_06514_),
    .S1(_06615_),
    .X(_06999_));
 sky130_fd_sc_hd__o221a_1 _12647_ (.A1(_06995_),
    .A2(_06998_),
    .B1(_06999_),
    .B2(_06824_),
    .C1(_06701_),
    .X(_07000_));
 sky130_fd_sc_hd__buf_12 _12648_ (.A(_06415_),
    .X(_07001_));
 sky130_fd_sc_hd__mux4_2 _12649_ (.A0(\fifo0.fifo_store[8][12] ),
    .A1(\fifo0.fifo_store[9][12] ),
    .A2(\fifo0.fifo_store[10][12] ),
    .A3(\fifo0.fifo_store[11][12] ),
    .S0(_07001_),
    .S1(_06691_),
    .X(_07002_));
 sky130_fd_sc_hd__mux4_1 _12650_ (.A0(\fifo0.fifo_store[12][12] ),
    .A1(\fifo0.fifo_store[13][12] ),
    .A2(\fifo0.fifo_store[14][12] ),
    .A3(\fifo0.fifo_store[15][12] ),
    .S0(_06513_),
    .S1(_06731_),
    .X(_07003_));
 sky130_fd_sc_hd__or2_1 _12651_ (.A(_06721_),
    .B(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__o211a_1 _12652_ (.A1(_06688_),
    .A2(_07002_),
    .B1(_07004_),
    .C1(_06686_),
    .X(_07005_));
 sky130_fd_sc_hd__mux4_1 _12653_ (.A0(\fifo0.fifo_store[24][12] ),
    .A1(\fifo0.fifo_store[25][12] ),
    .A2(\fifo0.fifo_store[26][12] ),
    .A3(\fifo0.fifo_store[27][12] ),
    .S0(_06415_),
    .S1(_06984_),
    .X(_07006_));
 sky130_fd_sc_hd__or2_1 _12654_ (.A(_06531_),
    .B(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__buf_12 _12655_ (.A(_06414_),
    .X(_07008_));
 sky130_fd_sc_hd__mux4_1 _12656_ (.A0(\fifo0.fifo_store[28][12] ),
    .A1(\fifo0.fifo_store[29][12] ),
    .A2(\fifo0.fifo_store[30][12] ),
    .A3(\fifo0.fifo_store[31][12] ),
    .S0(_07008_),
    .S1(_06725_),
    .X(_07009_));
 sky130_fd_sc_hd__o21a_1 _12657_ (.A1(_06709_),
    .A2(_07009_),
    .B1(_06713_),
    .X(_07010_));
 sky130_fd_sc_hd__mux4_1 _12658_ (.A0(\fifo0.fifo_store[16][12] ),
    .A1(\fifo0.fifo_store[17][12] ),
    .A2(\fifo0.fifo_store[18][12] ),
    .A3(\fifo0.fifo_store[19][12] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_07011_));
 sky130_fd_sc_hd__or2_1 _12659_ (.A(_06531_),
    .B(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__mux4_1 _12660_ (.A0(\fifo0.fifo_store[20][12] ),
    .A1(\fifo0.fifo_store[21][12] ),
    .A2(\fifo0.fifo_store[22][12] ),
    .A3(\fifo0.fifo_store[23][12] ),
    .S0(_07008_),
    .S1(_06695_),
    .X(_07013_));
 sky130_fd_sc_hd__o21a_1 _12661_ (.A1(_06709_),
    .A2(_07013_),
    .B1(_06444_),
    .X(_07014_));
 sky130_fd_sc_hd__a221o_1 _12662_ (.A1(_07007_),
    .A2(_07010_),
    .B1(_07012_),
    .B2(_07014_),
    .C1(_06743_),
    .X(_07015_));
 sky130_fd_sc_hd__o311a_4 _12663_ (.A1(_06966_),
    .A2(_07000_),
    .A3(_07005_),
    .B1(_06498_),
    .C1(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__buf_12 _12664_ (.A(_06486_),
    .X(_07017_));
 sky130_fd_sc_hd__or2_1 _12665_ (.A(_07017_),
    .B(\fifo0.fifo_store[52][12] ),
    .X(_07018_));
 sky130_fd_sc_hd__o211a_1 _12666_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[53][12] ),
    .B1(_07018_),
    .C1(_06699_),
    .X(_07019_));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(\fifo0.fifo_store[54][12] ),
    .A1(\fifo0.fifo_store[55][12] ),
    .S(_06469_),
    .X(_07020_));
 sky130_fd_sc_hd__a21o_1 _12668_ (.A1(_06996_),
    .A2(_07020_),
    .B1(_06721_),
    .X(_07021_));
 sky130_fd_sc_hd__buf_12 _12669_ (.A(_06513_),
    .X(_07022_));
 sky130_fd_sc_hd__mux4_1 _12670_ (.A0(\fifo0.fifo_store[48][12] ),
    .A1(\fifo0.fifo_store[49][12] ),
    .A2(\fifo0.fifo_store[50][12] ),
    .A3(\fifo0.fifo_store[51][12] ),
    .S0(_07022_),
    .S1(_06648_),
    .X(_07023_));
 sky130_fd_sc_hd__o221a_1 _12671_ (.A1(_07019_),
    .A2(_07021_),
    .B1(_07023_),
    .B2(_06824_),
    .C1(_06701_),
    .X(_07024_));
 sky130_fd_sc_hd__mux4_1 _12672_ (.A0(\fifo0.fifo_store[56][12] ),
    .A1(\fifo0.fifo_store[57][12] ),
    .A2(\fifo0.fifo_store[58][12] ),
    .A3(\fifo0.fifo_store[59][12] ),
    .S0(_06416_),
    .S1(_06971_),
    .X(_07025_));
 sky130_fd_sc_hd__mux4_1 _12673_ (.A0(\fifo0.fifo_store[60][12] ),
    .A1(\fifo0.fifo_store[61][12] ),
    .A2(\fifo0.fifo_store[62][12] ),
    .A3(\fifo0.fifo_store[63][12] ),
    .S0(_06617_),
    .S1(_06690_),
    .X(_07026_));
 sky130_fd_sc_hd__or2_1 _12674_ (.A(_06721_),
    .B(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__o211a_1 _12675_ (.A1(_06688_),
    .A2(_07025_),
    .B1(_07027_),
    .C1(_06686_),
    .X(_07028_));
 sky130_fd_sc_hd__mux4_1 _12676_ (.A0(\fifo0.fifo_store[40][12] ),
    .A1(\fifo0.fifo_store[41][12] ),
    .A2(\fifo0.fifo_store[42][12] ),
    .A3(\fifo0.fifo_store[43][12] ),
    .S0(_06617_),
    .S1(_06690_),
    .X(_07029_));
 sky130_fd_sc_hd__or2_1 _12677_ (.A(_06531_),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__mux4_2 _12678_ (.A0(\fifo0.fifo_store[44][12] ),
    .A1(\fifo0.fifo_store[45][12] ),
    .A2(\fifo0.fifo_store[46][12] ),
    .A3(\fifo0.fifo_store[47][12] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_07031_));
 sky130_fd_sc_hd__o21a_1 _12679_ (.A1(_06709_),
    .A2(_07031_),
    .B1(_06713_),
    .X(_07032_));
 sky130_fd_sc_hd__mux4_1 _12680_ (.A0(\fifo0.fifo_store[36][12] ),
    .A1(\fifo0.fifo_store[37][12] ),
    .A2(\fifo0.fifo_store[38][12] ),
    .A3(\fifo0.fifo_store[39][12] ),
    .S0(_06415_),
    .S1(_06984_),
    .X(_07033_));
 sky130_fd_sc_hd__or2_1 _12681_ (.A(_06721_),
    .B(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__mux4_1 _12682_ (.A0(\fifo0.fifo_store[32][12] ),
    .A1(\fifo0.fifo_store[33][12] ),
    .A2(\fifo0.fifo_store[34][12] ),
    .A3(\fifo0.fifo_store[35][12] ),
    .S0(_07008_),
    .S1(_06725_),
    .X(_07035_));
 sky130_fd_sc_hd__o21a_1 _12683_ (.A1(_06565_),
    .A2(_07035_),
    .B1(_06444_),
    .X(_07036_));
 sky130_fd_sc_hd__a221o_1 _12684_ (.A1(_07030_),
    .A2(_07032_),
    .B1(_07034_),
    .B2(_07036_),
    .C1(_06408_),
    .X(_07037_));
 sky130_fd_sc_hd__o311a_4 _12685_ (.A1(_06679_),
    .A2(_07024_),
    .A3(_07028_),
    .B1(_07037_),
    .C1(_06465_),
    .X(_07038_));
 sky130_fd_sc_hd__o31ai_1 _12686_ (.A1(_06992_),
    .A2(_07016_),
    .A3(_07038_),
    .B1(_06357_),
    .Y(_07039_));
 sky130_fd_sc_hd__o2bb2a_1 _12687_ (.A1_N(_06918_),
    .A2_N(_06938_),
    .B1(_06991_),
    .B2(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__a31o_1 _12688_ (.A1(_06377_),
    .A2(_06757_),
    .A3(_06786_),
    .B1(_06911_),
    .X(_07041_));
 sky130_fd_sc_hd__and2_1 _12689_ (.A(_06376_),
    .B(_06364_),
    .X(_07042_));
 sky130_fd_sc_hd__a21oi_1 _12690_ (.A1(_06382_),
    .A2(_06922_),
    .B1(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(_07041_),
    .A1(_07043_),
    .S(_06358_),
    .X(_07044_));
 sky130_fd_sc_hd__or2_1 _12692_ (.A(_06747_),
    .B(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__o21a_1 _12693_ (.A1(_06753_),
    .A2(_06927_),
    .B1(_06402_),
    .X(_07046_));
 sky130_fd_sc_hd__o211ai_1 _12694_ (.A1(_06392_),
    .A2(_06912_),
    .B1(_06786_),
    .C1(_06386_),
    .Y(_07047_));
 sky130_fd_sc_hd__o211a_1 _12695_ (.A1(_06922_),
    .A2(_07042_),
    .B1(_06923_),
    .C1(_06358_),
    .X(_07048_));
 sky130_fd_sc_hd__a211o_1 _12696_ (.A1(_07046_),
    .A2(_07047_),
    .B1(_07048_),
    .C1(_06769_),
    .X(_07049_));
 sky130_fd_sc_hd__a21oi_1 _12697_ (.A1(_06386_),
    .A2(_06753_),
    .B1(_06396_),
    .Y(_07050_));
 sky130_fd_sc_hd__a21o_1 _12698_ (.A1(_06396_),
    .A2(_06887_),
    .B1(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__o211a_1 _12699_ (.A1(_06398_),
    .A2(_06784_),
    .B1(_06761_),
    .C1(_06363_),
    .X(_07052_));
 sky130_fd_sc_hd__nor2_1 _12700_ (.A(_06902_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_06778_),
    .B(_06786_),
    .Y(_07054_));
 sky130_fd_sc_hd__a221o_1 _12702_ (.A1(_06359_),
    .A2(_07051_),
    .B1(_07053_),
    .B2(_07054_),
    .C1(_06747_),
    .X(_07055_));
 sky130_fd_sc_hd__xor2_2 _12703_ (.A(_06390_),
    .B(_06756_),
    .X(_07056_));
 sky130_fd_sc_hd__a21oi_2 _12704_ (.A1(_06748_),
    .A2(_06361_),
    .B1(_06395_),
    .Y(_07057_));
 sky130_fd_sc_hd__nand2_1 _12705_ (.A(_06398_),
    .B(_06761_),
    .Y(_07058_));
 sky130_fd_sc_hd__a221o_1 _12706_ (.A1(_06911_),
    .A2(_07056_),
    .B1(_07057_),
    .B2(_07058_),
    .C1(_06358_),
    .X(_07059_));
 sky130_fd_sc_hd__a211o_1 _12707_ (.A1(_06778_),
    .A2(_06779_),
    .B1(_07050_),
    .C1(_06402_),
    .X(_07060_));
 sky130_fd_sc_hd__a31oi_1 _12708_ (.A1(_06747_),
    .A2(_07059_),
    .A3(_07060_),
    .B1(_06405_),
    .Y(_07061_));
 sky130_fd_sc_hd__a32o_2 _12709_ (.A1(_06405_),
    .A2(_07045_),
    .A3(_07049_),
    .B1(_07055_),
    .B2(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__mux4_2 _12710_ (.A0(\fifo0.fifo_store[96][11] ),
    .A1(\fifo0.fifo_store[97][11] ),
    .A2(\fifo0.fifo_store[98][11] ),
    .A3(\fifo0.fifo_store[99][11] ),
    .S0(_06946_),
    .S1(_06648_),
    .X(_07063_));
 sky130_fd_sc_hd__mux4_1 _12711_ (.A0(\fifo0.fifo_store[100][11] ),
    .A1(\fifo0.fifo_store[101][11] ),
    .A2(\fifo0.fifo_store[102][11] ),
    .A3(\fifo0.fifo_store[103][11] ),
    .S0(_06946_),
    .S1(_06648_),
    .X(_07064_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(_07063_),
    .A1(_07064_),
    .S(_06656_),
    .X(_07065_));
 sky130_fd_sc_hd__buf_8 _12713_ (.A(_06565_),
    .X(_07066_));
 sky130_fd_sc_hd__buf_12 _12714_ (.A(_07008_),
    .X(_07067_));
 sky130_fd_sc_hd__mux4_1 _12715_ (.A0(\fifo0.fifo_store[104][11] ),
    .A1(\fifo0.fifo_store[105][11] ),
    .A2(\fifo0.fifo_store[106][11] ),
    .A3(\fifo0.fifo_store[107][11] ),
    .S0(_07067_),
    .S1(_06971_),
    .X(_07068_));
 sky130_fd_sc_hd__or2_1 _12716_ (.A(_07066_),
    .B(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__buf_8 _12717_ (.A(_06430_),
    .X(_07070_));
 sky130_fd_sc_hd__clkbuf_16 _12718_ (.A(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__buf_6 _12719_ (.A(_06470_),
    .X(_07072_));
 sky130_fd_sc_hd__buf_12 _12720_ (.A(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__mux4_1 _12721_ (.A0(\fifo0.fifo_store[108][11] ),
    .A1(\fifo0.fifo_store[109][11] ),
    .A2(\fifo0.fifo_store[110][11] ),
    .A3(\fifo0.fifo_store[111][11] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__o21a_1 _12722_ (.A1(_07071_),
    .A2(_07074_),
    .B1(_06686_),
    .X(_07075_));
 sky130_fd_sc_hd__a221o_1 _12723_ (.A1(_06939_),
    .A2(_07065_),
    .B1(_07069_),
    .B2(_07075_),
    .C1(_06966_),
    .X(_07076_));
 sky130_fd_sc_hd__buf_6 _12724_ (.A(_06412_),
    .X(_07077_));
 sky130_fd_sc_hd__or2_1 _12725_ (.A(_07077_),
    .B(\fifo0.fifo_store[119][11] ),
    .X(_07078_));
 sky130_fd_sc_hd__buf_12 _12726_ (.A(_06973_),
    .X(_07079_));
 sky130_fd_sc_hd__o21a_1 _12727_ (.A1(_07079_),
    .A2(\fifo0.fifo_store[118][11] ),
    .B1(_06996_),
    .X(_07080_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(\fifo0.fifo_store[116][11] ),
    .A1(\fifo0.fifo_store[117][11] ),
    .S(_06452_),
    .X(_07081_));
 sky130_fd_sc_hd__a221o_1 _12729_ (.A1(_07078_),
    .A2(_07080_),
    .B1(_07081_),
    .B2(_06954_),
    .C1(_06945_),
    .X(_07082_));
 sky130_fd_sc_hd__mux4_2 _12730_ (.A0(\fifo0.fifo_store[112][11] ),
    .A1(\fifo0.fifo_store[113][11] ),
    .A2(\fifo0.fifo_store[114][11] ),
    .A3(\fifo0.fifo_store[115][11] ),
    .S0(_07001_),
    .S1(_06691_),
    .X(_07083_));
 sky130_fd_sc_hd__or2_1 _12731_ (.A(_06688_),
    .B(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_16 _12732_ (.A(_06743_),
    .X(_07085_));
 sky130_fd_sc_hd__mux4_1 _12733_ (.A0(\fifo0.fifo_store[124][11] ),
    .A1(\fifo0.fifo_store[125][11] ),
    .A2(\fifo0.fifo_store[126][11] ),
    .A3(\fifo0.fifo_store[127][11] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_07086_));
 sky130_fd_sc_hd__mux4_1 _12734_ (.A0(\fifo0.fifo_store[120][11] ),
    .A1(\fifo0.fifo_store[121][11] ),
    .A2(\fifo0.fifo_store[122][11] ),
    .A3(\fifo0.fifo_store[123][11] ),
    .S0(_07008_),
    .S1(_06725_),
    .X(_07087_));
 sky130_fd_sc_hd__or2_1 _12735_ (.A(_06565_),
    .B(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__o211a_1 _12736_ (.A1(_07071_),
    .A2(_07086_),
    .B1(_07088_),
    .C1(_06686_),
    .X(_07089_));
 sky130_fd_sc_hd__a311o_1 _12737_ (.A1(_06939_),
    .A2(_07082_),
    .A3(_07084_),
    .B1(_07085_),
    .C1(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__mux4_1 _12738_ (.A0(\fifo0.fifo_store[76][11] ),
    .A1(\fifo0.fifo_store[77][11] ),
    .A2(\fifo0.fifo_store[78][11] ),
    .A3(\fifo0.fifo_store[79][11] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_07091_));
 sky130_fd_sc_hd__mux4_1 _12739_ (.A0(\fifo0.fifo_store[72][11] ),
    .A1(\fifo0.fifo_store[73][11] ),
    .A2(\fifo0.fifo_store[74][11] ),
    .A3(\fifo0.fifo_store[75][11] ),
    .S0(_06544_),
    .S1(_06695_),
    .X(_07092_));
 sky130_fd_sc_hd__or2_1 _12740_ (.A(_06565_),
    .B(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__clkbuf_16 _12741_ (.A(_06713_),
    .X(_07094_));
 sky130_fd_sc_hd__o211a_1 _12742_ (.A1(_07071_),
    .A2(_07091_),
    .B1(_07093_),
    .C1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__buf_12 _12743_ (.A(_06474_),
    .X(_07096_));
 sky130_fd_sc_hd__buf_12 _12744_ (.A(_06563_),
    .X(_07097_));
 sky130_fd_sc_hd__clkbuf_16 _12745_ (.A(_06470_),
    .X(_07098_));
 sky130_fd_sc_hd__buf_12 _12746_ (.A(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__mux4_2 _12747_ (.A0(\fifo0.fifo_store[64][11] ),
    .A1(\fifo0.fifo_store[65][11] ),
    .A2(\fifo0.fifo_store[66][11] ),
    .A3(\fifo0.fifo_store[67][11] ),
    .S0(_07097_),
    .S1(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__or2b_1 _12748_ (.A(\fifo0.fifo_store[71][11] ),
    .B_N(_07001_),
    .X(_07101_));
 sky130_fd_sc_hd__o21a_1 _12749_ (.A1(_07001_),
    .A2(\fifo0.fifo_store[70][11] ),
    .B1(_06504_),
    .X(_07102_));
 sky130_fd_sc_hd__mux2_1 _12750_ (.A0(\fifo0.fifo_store[68][11] ),
    .A1(\fifo0.fifo_store[69][11] ),
    .S(_06625_),
    .X(_07103_));
 sky130_fd_sc_hd__buf_8 _12751_ (.A(_06424_),
    .X(_07104_));
 sky130_fd_sc_hd__a221o_1 _12752_ (.A1(_07101_),
    .A2(_07102_),
    .B1(_07103_),
    .B2(_07104_),
    .C1(_07070_),
    .X(_07105_));
 sky130_fd_sc_hd__o211a_1 _12753_ (.A1(_07096_),
    .A2(_07100_),
    .B1(_07105_),
    .C1(_06445_),
    .X(_07106_));
 sky130_fd_sc_hd__buf_8 _12754_ (.A(_06444_),
    .X(_07107_));
 sky130_fd_sc_hd__mux4_1 _12755_ (.A0(\fifo0.fifo_store[80][11] ),
    .A1(\fifo0.fifo_store[81][11] ),
    .A2(\fifo0.fifo_store[82][11] ),
    .A3(\fifo0.fifo_store[83][11] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_07108_));
 sky130_fd_sc_hd__mux4_1 _12756_ (.A0(\fifo0.fifo_store[84][11] ),
    .A1(\fifo0.fifo_store[85][11] ),
    .A2(\fifo0.fifo_store[86][11] ),
    .A3(\fifo0.fifo_store[87][11] ),
    .S0(_06710_),
    .S1(_06711_),
    .X(_07109_));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(_07108_),
    .A1(_07109_),
    .S(_06730_),
    .X(_07110_));
 sky130_fd_sc_hd__buf_12 _12758_ (.A(_06470_),
    .X(_07111_));
 sky130_fd_sc_hd__mux4_1 _12759_ (.A0(\fifo0.fifo_store[88][11] ),
    .A1(\fifo0.fifo_store[89][11] ),
    .A2(\fifo0.fifo_store[90][11] ),
    .A3(\fifo0.fifo_store[91][11] ),
    .S0(_06563_),
    .S1(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__or2_1 _12760_ (.A(_06797_),
    .B(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__mux4_2 _12761_ (.A0(\fifo0.fifo_store[92][11] ),
    .A1(\fifo0.fifo_store[93][11] ),
    .A2(\fifo0.fifo_store[94][11] ),
    .A3(\fifo0.fifo_store[95][11] ),
    .S0(_06586_),
    .S1(_06471_),
    .X(_07114_));
 sky130_fd_sc_hd__o21a_1 _12762_ (.A1(_06431_),
    .A2(_07114_),
    .B1(_06713_),
    .X(_07115_));
 sky130_fd_sc_hd__a221o_1 _12763_ (.A1(_07107_),
    .A2(_07110_),
    .B1(_07113_),
    .B2(_07115_),
    .C1(_06539_),
    .X(_07116_));
 sky130_fd_sc_hd__o311a_1 _12764_ (.A1(_06966_),
    .A2(_07095_),
    .A3(_07106_),
    .B1(_07116_),
    .C1(_06498_),
    .X(_07117_));
 sky130_fd_sc_hd__a311oi_4 _12765_ (.A1(_06792_),
    .A2(_07076_),
    .A3(_07090_),
    .B1(_06965_),
    .C1(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__buf_8 _12766_ (.A(_06412_),
    .X(_07119_));
 sky130_fd_sc_hd__or2_1 _12767_ (.A(_06870_),
    .B(\fifo0.fifo_store[4][11] ),
    .X(_07120_));
 sky130_fd_sc_hd__o211a_1 _12768_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[5][11] ),
    .B1(_07120_),
    .C1(_07104_),
    .X(_07121_));
 sky130_fd_sc_hd__mux2_1 _12769_ (.A0(\fifo0.fifo_store[6][11] ),
    .A1(\fifo0.fifo_store[7][11] ),
    .S(_06600_),
    .X(_07122_));
 sky130_fd_sc_hd__a21o_1 _12770_ (.A1(_06454_),
    .A2(_07122_),
    .B1(_06709_),
    .X(_07123_));
 sky130_fd_sc_hd__mux4_1 _12771_ (.A0(\fifo0.fifo_store[0][11] ),
    .A1(\fifo0.fifo_store[1][11] ),
    .A2(\fifo0.fifo_store[2][11] ),
    .A3(\fifo0.fifo_store[3][11] ),
    .S0(_06416_),
    .S1(_06971_),
    .X(_07124_));
 sky130_fd_sc_hd__o221a_1 _12772_ (.A1(_07121_),
    .A2(_07123_),
    .B1(_07124_),
    .B2(_07066_),
    .C1(_07107_),
    .X(_07125_));
 sky130_fd_sc_hd__mux4_2 _12773_ (.A0(\fifo0.fifo_store[8][11] ),
    .A1(\fifo0.fifo_store[9][11] ),
    .A2(\fifo0.fifo_store[10][11] ),
    .A3(\fifo0.fifo_store[11][11] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_07126_));
 sky130_fd_sc_hd__mux4_1 _12774_ (.A0(\fifo0.fifo_store[12][11] ),
    .A1(\fifo0.fifo_store[13][11] ),
    .A2(\fifo0.fifo_store[14][11] ),
    .A3(\fifo0.fifo_store[15][11] ),
    .S0(_06544_),
    .S1(_06695_),
    .X(_07127_));
 sky130_fd_sc_hd__or2_1 _12775_ (.A(_06709_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__o211a_1 _12776_ (.A1(_07096_),
    .A2(_07126_),
    .B1(_07128_),
    .C1(_07094_),
    .X(_07129_));
 sky130_fd_sc_hd__mux4_1 _12777_ (.A0(\fifo0.fifo_store[24][11] ),
    .A1(\fifo0.fifo_store[25][11] ),
    .A2(\fifo0.fifo_store[26][11] ),
    .A3(\fifo0.fifo_store[27][11] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_07130_));
 sky130_fd_sc_hd__or2_1 _12778_ (.A(_06474_),
    .B(_07130_),
    .X(_07131_));
 sky130_fd_sc_hd__buf_12 _12779_ (.A(_06430_),
    .X(_07132_));
 sky130_fd_sc_hd__mux4_1 _12780_ (.A0(\fifo0.fifo_store[28][11] ),
    .A1(\fifo0.fifo_store[29][11] ),
    .A2(\fifo0.fifo_store[30][11] ),
    .A3(\fifo0.fifo_store[31][11] ),
    .S0(_06434_),
    .S1(_07098_),
    .X(_07133_));
 sky130_fd_sc_hd__o21a_1 _12781_ (.A1(_07132_),
    .A2(_07133_),
    .B1(_06713_),
    .X(_07134_));
 sky130_fd_sc_hd__mux4_1 _12782_ (.A0(\fifo0.fifo_store[16][11] ),
    .A1(\fifo0.fifo_store[17][11] ),
    .A2(\fifo0.fifo_store[18][11] ),
    .A3(\fifo0.fifo_store[19][11] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_07135_));
 sky130_fd_sc_hd__or2_1 _12783_ (.A(_06797_),
    .B(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__mux4_2 _12784_ (.A0(\fifo0.fifo_store[20][11] ),
    .A1(\fifo0.fifo_store[21][11] ),
    .A2(\fifo0.fifo_store[22][11] ),
    .A3(\fifo0.fifo_store[23][11] ),
    .S0(_06586_),
    .S1(_06471_),
    .X(_07137_));
 sky130_fd_sc_hd__o21a_1 _12785_ (.A1(_06431_),
    .A2(_07137_),
    .B1(_06444_),
    .X(_07138_));
 sky130_fd_sc_hd__a221o_1 _12786_ (.A1(_07131_),
    .A2(_07134_),
    .B1(_07136_),
    .B2(_07138_),
    .C1(_06539_),
    .X(_07139_));
 sky130_fd_sc_hd__o311a_4 _12787_ (.A1(_06966_),
    .A2(_07125_),
    .A3(_07129_),
    .B1(_06498_),
    .C1(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__or2_1 _12788_ (.A(_06549_),
    .B(\fifo0.fifo_store[52][11] ),
    .X(_07141_));
 sky130_fd_sc_hd__o211a_1 _12789_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[53][11] ),
    .B1(_07141_),
    .C1(_07104_),
    .X(_07142_));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(\fifo0.fifo_store[54][11] ),
    .A1(\fifo0.fifo_store[55][11] ),
    .S(_06569_),
    .X(_07143_));
 sky130_fd_sc_hd__a21o_1 _12791_ (.A1(_06454_),
    .A2(_07143_),
    .B1(_06709_),
    .X(_07144_));
 sky130_fd_sc_hd__mux4_1 _12792_ (.A0(\fifo0.fifo_store[48][11] ),
    .A1(\fifo0.fifo_store[49][11] ),
    .A2(\fifo0.fifo_store[50][11] ),
    .A3(\fifo0.fifo_store[51][11] ),
    .S0(_07067_),
    .S1(_06971_),
    .X(_07145_));
 sky130_fd_sc_hd__o221a_1 _12793_ (.A1(_07142_),
    .A2(_07144_),
    .B1(_07145_),
    .B2(_07066_),
    .C1(_07107_),
    .X(_07146_));
 sky130_fd_sc_hd__mux4_1 _12794_ (.A0(\fifo0.fifo_store[56][11] ),
    .A1(\fifo0.fifo_store[57][11] ),
    .A2(\fifo0.fifo_store[58][11] ),
    .A3(\fifo0.fifo_store[59][11] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_07147_));
 sky130_fd_sc_hd__mux4_1 _12795_ (.A0(\fifo0.fifo_store[60][11] ),
    .A1(\fifo0.fifo_store[61][11] ),
    .A2(\fifo0.fifo_store[62][11] ),
    .A3(\fifo0.fifo_store[63][11] ),
    .S0(_06507_),
    .S1(_07072_),
    .X(_07148_));
 sky130_fd_sc_hd__or2_1 _12796_ (.A(_07070_),
    .B(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__o211a_1 _12797_ (.A1(_07096_),
    .A2(_07147_),
    .B1(_07149_),
    .C1(_07094_),
    .X(_07150_));
 sky130_fd_sc_hd__mux4_1 _12798_ (.A0(\fifo0.fifo_store[40][11] ),
    .A1(\fifo0.fifo_store[41][11] ),
    .A2(\fifo0.fifo_store[42][11] ),
    .A3(\fifo0.fifo_store[43][11] ),
    .S0(_06507_),
    .S1(_06975_),
    .X(_07151_));
 sky130_fd_sc_hd__or2_1 _12799_ (.A(_06474_),
    .B(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__mux4_1 _12800_ (.A0(\fifo0.fifo_store[44][11] ),
    .A1(\fifo0.fifo_store[45][11] ),
    .A2(\fifo0.fifo_store[46][11] ),
    .A3(\fifo0.fifo_store[47][11] ),
    .S0(_06563_),
    .S1(_07111_),
    .X(_07153_));
 sky130_fd_sc_hd__o21a_1 _12801_ (.A1(_07132_),
    .A2(_07153_),
    .B1(_06713_),
    .X(_07154_));
 sky130_fd_sc_hd__mux4_1 _12802_ (.A0(\fifo0.fifo_store[36][11] ),
    .A1(\fifo0.fifo_store[37][11] ),
    .A2(\fifo0.fifo_store[38][11] ),
    .A3(\fifo0.fifo_store[39][11] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_07155_));
 sky130_fd_sc_hd__or2_1 _12803_ (.A(_07070_),
    .B(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__mux4_1 _12804_ (.A0(\fifo0.fifo_store[32][11] ),
    .A1(\fifo0.fifo_store[33][11] ),
    .A2(\fifo0.fifo_store[34][11] ),
    .A3(\fifo0.fifo_store[35][11] ),
    .S0(_06434_),
    .S1(_06561_),
    .X(_07157_));
 sky130_fd_sc_hd__o21a_1 _12805_ (.A1(_06441_),
    .A2(_07157_),
    .B1(_06444_),
    .X(_07158_));
 sky130_fd_sc_hd__a221o_1 _12806_ (.A1(_07152_),
    .A2(_07154_),
    .B1(_07156_),
    .B2(_07158_),
    .C1(_06408_),
    .X(_07159_));
 sky130_fd_sc_hd__o311a_4 _12807_ (.A1(_07085_),
    .A2(_07146_),
    .A3(_07150_),
    .B1(_07159_),
    .C1(_06465_),
    .X(_07160_));
 sky130_fd_sc_hd__o31ai_2 _12808_ (.A1(_06992_),
    .A2(_07140_),
    .A3(_07160_),
    .B1(_06357_),
    .Y(_07161_));
 sky130_fd_sc_hd__o22a_1 _12809_ (.A1(_06611_),
    .A2(_07062_),
    .B1(_07118_),
    .B2(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__clkinv_2 _12810_ (.A(net30),
    .Y(_07163_));
 sky130_fd_sc_hd__clkbuf_4 _12811_ (.A(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__inv_2 _12812_ (.A(net31),
    .Y(_07165_));
 sky130_fd_sc_hd__mux4_1 _12813_ (.A0(_06791_),
    .A1(_06917_),
    .A2(_07040_),
    .A3(_07162_),
    .S0(_07164_),
    .S1(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__nand2_2 _12814_ (.A(_06407_),
    .B(_06607_),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_1 _12815_ (.A(net32),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__o21a_1 _12816_ (.A1(net32),
    .A2(_07166_),
    .B1(_07168_),
    .X(_07169_));
 sky130_fd_sc_hd__inv_2 _12817_ (.A(net33),
    .Y(_07170_));
 sky130_fd_sc_hd__nor2_2 _12818_ (.A(net31),
    .B(net32),
    .Y(_07171_));
 sky130_fd_sc_hd__and3_1 _12819_ (.A(_07164_),
    .B(_07170_),
    .C(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__buf_2 _12820_ (.A(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__a21oi_1 _12821_ (.A1(_06354_),
    .A2(_07167_),
    .B1(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__o21ai_1 _12822_ (.A1(_06354_),
    .A2(_07169_),
    .B1(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_07173_),
    .A2(_07162_),
    .B1(_06356_),
    .Y(_07176_));
 sky130_fd_sc_hd__and2_1 _12824_ (.A(_07175_),
    .B(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__nor2_1 _12825_ (.A(\dsmod0.accu1[11] ),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__and3_1 _12826_ (.A(\dsmod0.accu1[11] ),
    .B(_07175_),
    .C(_07176_),
    .X(_07179_));
 sky130_fd_sc_hd__or2_1 _12827_ (.A(_07178_),
    .B(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__or4_1 _12828_ (.A(net31),
    .B(_06353_),
    .C(_06354_),
    .D(net32),
    .X(_07181_));
 sky130_fd_sc_hd__clkbuf_2 _12829_ (.A(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__a32o_1 _12830_ (.A1(_06396_),
    .A2(_06897_),
    .A3(_06766_),
    .B1(_07058_),
    .B2(_07057_),
    .X(_07183_));
 sky130_fd_sc_hd__nor3_1 _12831_ (.A(_06362_),
    .B(_06391_),
    .C(_06380_),
    .Y(_07184_));
 sky130_fd_sc_hd__a211o_1 _12832_ (.A1(_06363_),
    .A2(_07056_),
    .B1(_07184_),
    .C1(_06358_),
    .X(_07185_));
 sky130_fd_sc_hd__o211a_1 _12833_ (.A1(_06402_),
    .A2(_07183_),
    .B1(_07185_),
    .C1(_06405_),
    .X(_07186_));
 sky130_fd_sc_hd__o211a_1 _12834_ (.A1(_06886_),
    .A2(_06367_),
    .B1(_06910_),
    .C1(_07054_),
    .X(_07187_));
 sky130_fd_sc_hd__or3b_1 _12835_ (.A(_07057_),
    .B(_06374_),
    .C_N(_06934_),
    .X(_07188_));
 sky130_fd_sc_hd__nand2_1 _12836_ (.A(_06919_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__or3_1 _12837_ (.A(_07186_),
    .B(_07187_),
    .C(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__o21ai_1 _12838_ (.A1(_06886_),
    .A2(_06367_),
    .B1(_06397_),
    .Y(_07191_));
 sky130_fd_sc_hd__o211a_1 _12839_ (.A1(_06753_),
    .A2(_06927_),
    .B1(_06910_),
    .C1(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__nor2_1 _12840_ (.A(\sinegen0.read_ptr[5] ),
    .B(_06373_),
    .Y(_07193_));
 sky130_fd_sc_hd__o211a_1 _12841_ (.A1(_06392_),
    .A2(_06912_),
    .B1(_07193_),
    .C1(_06772_),
    .X(_07194_));
 sky130_fd_sc_hd__or3b_1 _12842_ (.A(_06362_),
    .B(_06391_),
    .C_N(_06761_),
    .X(_07195_));
 sky130_fd_sc_hd__o2111a_1 _12843_ (.A1(_06393_),
    .A2(_06923_),
    .B1(_07195_),
    .C1(_06401_),
    .D1(_06404_),
    .X(_07196_));
 sky130_fd_sc_hd__or4_1 _12844_ (.A(\sinegen0.read_ptr[6] ),
    .B(_07192_),
    .C(_07194_),
    .D(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__nand2_1 _12845_ (.A(_06404_),
    .B(_06902_),
    .Y(_07198_));
 sky130_fd_sc_hd__a221o_1 _12846_ (.A1(_06891_),
    .A2(_06751_),
    .B1(_07058_),
    .B2(_07057_),
    .C1(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__or2b_1 _12847_ (.A(_07197_),
    .B_N(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__a21o_1 _12848_ (.A1(_07190_),
    .A2(_07200_),
    .B1(_06606_),
    .X(_07201_));
 sky130_fd_sc_hd__buf_8 _12849_ (.A(_06804_),
    .X(_07202_));
 sky130_fd_sc_hd__buf_8 _12850_ (.A(_07096_),
    .X(_07203_));
 sky130_fd_sc_hd__buf_8 _12851_ (.A(_07067_),
    .X(_07204_));
 sky130_fd_sc_hd__buf_12 _12852_ (.A(_06648_),
    .X(_07205_));
 sky130_fd_sc_hd__mux4_1 _12853_ (.A0(\fifo0.fifo_store[48][10] ),
    .A1(\fifo0.fifo_store[49][10] ),
    .A2(\fifo0.fifo_store[50][10] ),
    .A3(\fifo0.fifo_store[51][10] ),
    .S0(_07204_),
    .S1(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__buf_8 _12854_ (.A(_06954_),
    .X(_07207_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(\fifo0.fifo_store[52][10] ),
    .A1(\fifo0.fifo_store[53][10] ),
    .S(_07079_),
    .X(_07208_));
 sky130_fd_sc_hd__buf_12 _12856_ (.A(_06615_),
    .X(_07209_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(\fifo0.fifo_store[54][10] ),
    .A1(\fifo0.fifo_store[55][10] ),
    .S(_07022_),
    .X(_07210_));
 sky130_fd_sc_hd__a21o_1 _12858_ (.A1(_07209_),
    .A2(_07210_),
    .B1(_06502_),
    .X(_07211_));
 sky130_fd_sc_hd__a21o_1 _12859_ (.A1(_07207_),
    .A2(_07208_),
    .B1(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__o211ai_1 _12860_ (.A1(_07203_),
    .A2(_07206_),
    .B1(_07212_),
    .C1(_06939_),
    .Y(_07213_));
 sky130_fd_sc_hd__mux4_1 _12861_ (.A0(\fifo0.fifo_store[56][10] ),
    .A1(\fifo0.fifo_store[57][10] ),
    .A2(\fifo0.fifo_store[58][10] ),
    .A3(\fifo0.fifo_store[59][10] ),
    .S0(_07204_),
    .S1(_07205_),
    .X(_07214_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(\fifo0.fifo_store[60][10] ),
    .A1(\fifo0.fifo_store[61][10] ),
    .S(_07079_),
    .X(_07215_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(\fifo0.fifo_store[62][10] ),
    .A1(\fifo0.fifo_store[63][10] ),
    .S(_06959_),
    .X(_07216_));
 sky130_fd_sc_hd__a21o_1 _12864_ (.A1(_07209_),
    .A2(_07216_),
    .B1(_06502_),
    .X(_07217_));
 sky130_fd_sc_hd__a21o_1 _12865_ (.A1(_06954_),
    .A2(_07215_),
    .B1(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__buf_6 _12866_ (.A(_06461_),
    .X(_07219_));
 sky130_fd_sc_hd__buf_8 _12867_ (.A(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__o211ai_1 _12868_ (.A1(_07203_),
    .A2(_07214_),
    .B1(_07218_),
    .C1(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__mux4_1 _12869_ (.A0(\fifo0.fifo_store[40][10] ),
    .A1(\fifo0.fifo_store[41][10] ),
    .A2(\fifo0.fifo_store[42][10] ),
    .A3(\fifo0.fifo_store[43][10] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_07222_));
 sky130_fd_sc_hd__or2_1 _12870_ (.A(_07096_),
    .B(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__mux4_1 _12871_ (.A0(\fifo0.fifo_store[44][10] ),
    .A1(\fifo0.fifo_store[45][10] ),
    .A2(\fifo0.fifo_store[46][10] ),
    .A3(\fifo0.fifo_store[47][10] ),
    .S0(_07097_),
    .S1(_07099_),
    .X(_07224_));
 sky130_fd_sc_hd__o21a_1 _12872_ (.A1(_07071_),
    .A2(_07224_),
    .B1(_07094_),
    .X(_07225_));
 sky130_fd_sc_hd__buf_8 _12873_ (.A(_06412_),
    .X(_07226_));
 sky130_fd_sc_hd__buf_12 _12874_ (.A(_06717_),
    .X(_07227_));
 sky130_fd_sc_hd__or2_1 _12875_ (.A(_07227_),
    .B(\fifo0.fifo_store[36][10] ),
    .X(_07228_));
 sky130_fd_sc_hd__o211a_1 _12876_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[37][10] ),
    .B1(_07228_),
    .C1(_07104_),
    .X(_07229_));
 sky130_fd_sc_hd__mux2_1 _12877_ (.A0(\fifo0.fifo_store[38][10] ),
    .A1(\fifo0.fifo_store[39][10] ),
    .S(_07017_),
    .X(_07230_));
 sky130_fd_sc_hd__a21o_1 _12878_ (.A1(_06556_),
    .A2(_07230_),
    .B1(_07070_),
    .X(_07231_));
 sky130_fd_sc_hd__mux4_2 _12879_ (.A0(\fifo0.fifo_store[32][10] ),
    .A1(\fifo0.fifo_store[33][10] ),
    .A2(\fifo0.fifo_store[34][10] ),
    .A3(\fifo0.fifo_store[35][10] ),
    .S0(_06545_),
    .S1(_07073_),
    .X(_07232_));
 sky130_fd_sc_hd__o221a_1 _12880_ (.A1(_07229_),
    .A2(_07231_),
    .B1(_07232_),
    .B2(_07066_),
    .C1(_07107_),
    .X(_07233_));
 sky130_fd_sc_hd__a211oi_2 _12881_ (.A1(_07223_),
    .A2(_07225_),
    .B1(_07233_),
    .C1(_06409_),
    .Y(_07234_));
 sky130_fd_sc_hd__a311o_4 _12882_ (.A1(_07202_),
    .A2(_07213_),
    .A3(_07221_),
    .B1(_06575_),
    .C1(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__mux4_1 _12883_ (.A0(\fifo0.fifo_store[20][10] ),
    .A1(\fifo0.fifo_store[21][10] ),
    .A2(\fifo0.fifo_store[22][10] ),
    .A3(\fifo0.fifo_store[23][10] ),
    .S0(_06545_),
    .S1(_07073_),
    .X(_07236_));
 sky130_fd_sc_hd__nor2_1 _12884_ (.A(_06945_),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__mux4_2 _12885_ (.A0(\fifo0.fifo_store[16][10] ),
    .A1(\fifo0.fifo_store[17][10] ),
    .A2(\fifo0.fifo_store[18][10] ),
    .A3(\fifo0.fifo_store[19][10] ),
    .S0(_06689_),
    .S1(_06691_),
    .X(_07238_));
 sky130_fd_sc_hd__o21ai_1 _12886_ (.A1(_06688_),
    .A2(_07238_),
    .B1(_06701_),
    .Y(_07239_));
 sky130_fd_sc_hd__mux4_2 _12887_ (.A0(\fifo0.fifo_store[24][10] ),
    .A1(\fifo0.fifo_store[25][10] ),
    .A2(\fifo0.fifo_store[26][10] ),
    .A3(\fifo0.fifo_store[27][10] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_07240_));
 sky130_fd_sc_hd__nor2_1 _12888_ (.A(_07066_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__mux4_1 _12889_ (.A0(\fifo0.fifo_store[28][10] ),
    .A1(\fifo0.fifo_store[29][10] ),
    .A2(\fifo0.fifo_store[30][10] ),
    .A3(\fifo0.fifo_store[31][10] ),
    .S0(_06416_),
    .S1(_06691_),
    .X(_07242_));
 sky130_fd_sc_hd__o21ai_1 _12890_ (.A1(_06945_),
    .A2(_07242_),
    .B1(_06686_),
    .Y(_07243_));
 sky130_fd_sc_hd__o221a_1 _12891_ (.A1(_07237_),
    .A2(_07239_),
    .B1(_07241_),
    .B2(_07243_),
    .C1(_06804_),
    .X(_07244_));
 sky130_fd_sc_hd__mux4_1 _12892_ (.A0(\fifo0.fifo_store[12][10] ),
    .A1(\fifo0.fifo_store[13][10] ),
    .A2(\fifo0.fifo_store[14][10] ),
    .A3(\fifo0.fifo_store[15][10] ),
    .S0(_06795_),
    .S1(_06504_),
    .X(_07245_));
 sky130_fd_sc_hd__or2_1 _12893_ (.A(_06502_),
    .B(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__mux4_1 _12894_ (.A0(\fifo0.fifo_store[8][10] ),
    .A1(\fifo0.fifo_store[9][10] ),
    .A2(\fifo0.fifo_store[10][10] ),
    .A3(\fifo0.fifo_store[11][10] ),
    .S0(_06479_),
    .S1(_06811_),
    .X(_07247_));
 sky130_fd_sc_hd__o21a_1 _12895_ (.A1(_06599_),
    .A2(_07247_),
    .B1(_06571_),
    .X(_07248_));
 sky130_fd_sc_hd__mux4_1 _12896_ (.A0(\fifo0.fifo_store[4][10] ),
    .A1(\fifo0.fifo_store[5][10] ),
    .A2(\fifo0.fifo_store[6][10] ),
    .A3(\fifo0.fifo_store[7][10] ),
    .S0(_06591_),
    .S1(_06592_),
    .X(_07249_));
 sky130_fd_sc_hd__mux4_1 _12897_ (.A0(\fifo0.fifo_store[0][10] ),
    .A1(\fifo0.fifo_store[1][10] ),
    .A2(\fifo0.fifo_store[2][10] ),
    .A3(\fifo0.fifo_store[3][10] ),
    .S0(_06977_),
    .S1(_06592_),
    .X(_07250_));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(_07249_),
    .A1(_07250_),
    .S(_07070_),
    .X(_07251_));
 sky130_fd_sc_hd__a221o_1 _12899_ (.A1(_07246_),
    .A2(_07248_),
    .B1(_07251_),
    .B2(_06552_),
    .C1(_06589_),
    .X(_07252_));
 sky130_fd_sc_hd__or3b_4 _12900_ (.A(_06465_),
    .B(_07244_),
    .C_N(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__mux4_1 _12901_ (.A0(\fifo0.fifo_store[88][10] ),
    .A1(\fifo0.fifo_store[89][10] ),
    .A2(\fifo0.fifo_store[90][10] ),
    .A3(\fifo0.fifo_store[91][10] ),
    .S0(_06545_),
    .S1(_07073_),
    .X(_07254_));
 sky130_fd_sc_hd__or2_1 _12902_ (.A(_06946_),
    .B(\fifo0.fifo_store[92][10] ),
    .X(_07255_));
 sky130_fd_sc_hd__o211a_1 _12903_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[93][10] ),
    .B1(_07255_),
    .C1(_06516_),
    .X(_07256_));
 sky130_fd_sc_hd__buf_12 _12904_ (.A(_06511_),
    .X(_07257_));
 sky130_fd_sc_hd__mux2_1 _12905_ (.A0(\fifo0.fifo_store[94][10] ),
    .A1(\fifo0.fifo_store[95][10] ),
    .S(_06549_),
    .X(_07258_));
 sky130_fd_sc_hd__a21o_1 _12906_ (.A1(_07257_),
    .A2(_07258_),
    .B1(_06431_),
    .X(_07259_));
 sky130_fd_sc_hd__o22a_1 _12907_ (.A1(_07066_),
    .A2(_07254_),
    .B1(_07256_),
    .B2(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__or2_1 _12908_ (.A(_06427_),
    .B(\fifo0.fifo_store[86][10] ),
    .X(_07261_));
 sky130_fd_sc_hd__o211a_1 _12909_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[87][10] ),
    .B1(_07261_),
    .C1(_06454_),
    .X(_07262_));
 sky130_fd_sc_hd__buf_12 _12910_ (.A(_06478_),
    .X(_07263_));
 sky130_fd_sc_hd__mux2_1 _12911_ (.A0(\fifo0.fifo_store[84][10] ),
    .A1(\fifo0.fifo_store[85][10] ),
    .S(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__a21o_1 _12912_ (.A1(_07104_),
    .A2(_07264_),
    .B1(_07070_),
    .X(_07265_));
 sky130_fd_sc_hd__mux4_1 _12913_ (.A0(\fifo0.fifo_store[80][10] ),
    .A1(\fifo0.fifo_store[81][10] ),
    .A2(\fifo0.fifo_store[82][10] ),
    .A3(\fifo0.fifo_store[83][10] ),
    .S0(_06545_),
    .S1(_06971_),
    .X(_07266_));
 sky130_fd_sc_hd__o221a_1 _12914_ (.A1(_07262_),
    .A2(_07265_),
    .B1(_07266_),
    .B2(_07066_),
    .C1(_07107_),
    .X(_07267_));
 sky130_fd_sc_hd__a211oi_1 _12915_ (.A1(_07220_),
    .A2(_07260_),
    .B1(_07267_),
    .C1(_07085_),
    .Y(_07268_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(\fifo0.fifo_store[76][10] ),
    .A1(\fifo0.fifo_store[77][10] ),
    .S(_06959_),
    .X(_07269_));
 sky130_fd_sc_hd__nand2_1 _12917_ (.A(_06954_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(\fifo0.fifo_store[78][10] ),
    .A1(\fifo0.fifo_store[79][10] ),
    .S(_06959_),
    .X(_07271_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(_07209_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__mux4_1 _12920_ (.A0(\fifo0.fifo_store[72][10] ),
    .A1(\fifo0.fifo_store[73][10] ),
    .A2(\fifo0.fifo_store[74][10] ),
    .A3(\fifo0.fifo_store[75][10] ),
    .S0(_06563_),
    .S1(_06561_),
    .X(_07273_));
 sky130_fd_sc_hd__o21ai_1 _12921_ (.A1(_06797_),
    .A2(_07273_),
    .B1(_06462_),
    .Y(_07274_));
 sky130_fd_sc_hd__a31o_1 _12922_ (.A1(_06688_),
    .A2(_07270_),
    .A3(_07272_),
    .B1(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__or2_1 _12923_ (.A(_06427_),
    .B(\fifo0.fifo_store[68][10] ),
    .X(_07276_));
 sky130_fd_sc_hd__o211a_1 _12924_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[69][10] ),
    .B1(_07276_),
    .C1(_07104_),
    .X(_07277_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(\fifo0.fifo_store[70][10] ),
    .A1(\fifo0.fifo_store[71][10] ),
    .S(_06487_),
    .X(_07278_));
 sky130_fd_sc_hd__a21o_1 _12926_ (.A1(_06556_),
    .A2(_07278_),
    .B1(_07070_),
    .X(_07279_));
 sky130_fd_sc_hd__mux4_2 _12927_ (.A0(\fifo0.fifo_store[64][10] ),
    .A1(\fifo0.fifo_store[65][10] ),
    .A2(\fifo0.fifo_store[66][10] ),
    .A3(\fifo0.fifo_store[67][10] ),
    .S0(_07067_),
    .S1(_06971_),
    .X(_07280_));
 sky130_fd_sc_hd__o221ai_1 _12928_ (.A1(_07277_),
    .A2(_07279_),
    .B1(_07280_),
    .B2(_07096_),
    .C1(_07107_),
    .Y(_07281_));
 sky130_fd_sc_hd__a31o_1 _12929_ (.A1(_06679_),
    .A2(_07275_),
    .A3(_07281_),
    .B1(_00005_),
    .X(_07282_));
 sky130_fd_sc_hd__mux4_2 _12930_ (.A0(\fifo0.fifo_store[112][10] ),
    .A1(\fifo0.fifo_store[113][10] ),
    .A2(\fifo0.fifo_store[114][10] ),
    .A3(\fifo0.fifo_store[115][10] ),
    .S0(_06801_),
    .S1(_06421_),
    .X(_07283_));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(\fifo0.fifo_store[116][10] ),
    .A1(\fifo0.fifo_store[117][10] ),
    .S(_06801_),
    .X(_07284_));
 sky130_fd_sc_hd__nand2_1 _12932_ (.A(_06425_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(\fifo0.fifo_store[118][10] ),
    .A1(\fifo0.fifo_store[119][10] ),
    .S(_06479_),
    .X(_07286_));
 sky130_fd_sc_hd__a21oi_1 _12934_ (.A1(_06556_),
    .A2(_07286_),
    .B1(_07070_),
    .Y(_07287_));
 sky130_fd_sc_hd__a2bb2o_1 _12935_ (.A1_N(_06624_),
    .A2_N(_07283_),
    .B1(_07285_),
    .B2(_07287_),
    .X(_07288_));
 sky130_fd_sc_hd__mux4_2 _12936_ (.A0(\fifo0.fifo_store[120][10] ),
    .A1(\fifo0.fifo_store[121][10] ),
    .A2(\fifo0.fifo_store[122][10] ),
    .A3(\fifo0.fifo_store[123][10] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_07289_));
 sky130_fd_sc_hd__nor2_1 _12937_ (.A(_06449_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(\fifo0.fifo_store[124][10] ),
    .A1(\fifo0.fifo_store[125][10] ),
    .S(_07227_),
    .X(_07291_));
 sky130_fd_sc_hd__nand2_1 _12939_ (.A(_06954_),
    .B(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(\fifo0.fifo_store[126][10] ),
    .A1(\fifo0.fifo_store[127][10] ),
    .S(_07227_),
    .X(_07293_));
 sky130_fd_sc_hd__nand2_1 _12941_ (.A(_07209_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__a31o_1 _12942_ (.A1(_06824_),
    .A2(_07292_),
    .A3(_07294_),
    .B1(_06735_),
    .X(_07295_));
 sky130_fd_sc_hd__o221a_1 _12943_ (.A1(_07220_),
    .A2(_07288_),
    .B1(_07290_),
    .B2(_07295_),
    .C1(_06966_),
    .X(_07296_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(\fifo0.fifo_store[110][10] ),
    .A1(\fifo0.fifo_store[111][10] ),
    .S(_06946_),
    .X(_07297_));
 sky130_fd_sc_hd__nand2_1 _12945_ (.A(_07205_),
    .B(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(\fifo0.fifo_store[108][10] ),
    .A1(\fifo0.fifo_store[109][10] ),
    .S(_06658_),
    .X(_07299_));
 sky130_fd_sc_hd__a21oi_1 _12947_ (.A1(_06425_),
    .A2(_07299_),
    .B1(_06431_),
    .Y(_07300_));
 sky130_fd_sc_hd__mux4_1 _12948_ (.A0(\fifo0.fifo_store[104][10] ),
    .A1(\fifo0.fifo_store[105][10] ),
    .A2(\fifo0.fifo_store[106][10] ),
    .A3(\fifo0.fifo_store[107][10] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_07301_));
 sky130_fd_sc_hd__nor2_1 _12949_ (.A(_06519_),
    .B(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__a211o_1 _12950_ (.A1(_07298_),
    .A2(_07300_),
    .B1(_06735_),
    .C1(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__or2_1 _12951_ (.A(_06514_),
    .B(\fifo0.fifo_store[102][10] ),
    .X(_07304_));
 sky130_fd_sc_hd__o211a_1 _12952_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[103][10] ),
    .B1(_07304_),
    .C1(_06556_),
    .X(_07305_));
 sky130_fd_sc_hd__mux2_1 _12953_ (.A0(\fifo0.fifo_store[100][10] ),
    .A1(\fifo0.fifo_store[101][10] ),
    .S(_06848_),
    .X(_07306_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_06516_),
    .A2(_07306_),
    .B1(_07132_),
    .X(_07307_));
 sky130_fd_sc_hd__mux4_2 _12955_ (.A0(\fifo0.fifo_store[96][10] ),
    .A1(\fifo0.fifo_store[97][10] ),
    .A2(\fifo0.fifo_store[98][10] ),
    .A3(\fifo0.fifo_store[99][10] ),
    .S0(_06545_),
    .S1(_07073_),
    .X(_07308_));
 sky130_fd_sc_hd__o221ai_1 _12956_ (.A1(_07305_),
    .A2(_07307_),
    .B1(_07308_),
    .B2(_07096_),
    .C1(_07107_),
    .Y(_07309_));
 sky130_fd_sc_hd__a31o_1 _12957_ (.A1(_06679_),
    .A2(_07303_),
    .A3(_07309_),
    .B1(_06677_),
    .X(_07310_));
 sky130_fd_sc_hd__o221a_4 _12958_ (.A1(_07268_),
    .A2(_07282_),
    .B1(_07296_),
    .B2(_07310_),
    .C1(_06992_),
    .X(_07311_));
 sky130_fd_sc_hd__a311o_2 _12959_ (.A1(_06965_),
    .A2(_07235_),
    .A3(_07253_),
    .B1(_07311_),
    .C1(_06918_),
    .X(_07312_));
 sky130_fd_sc_hd__nand2_1 _12960_ (.A(_07201_),
    .B(_07312_),
    .Y(_07313_));
 sky130_fd_sc_hd__buf_2 _12961_ (.A(_07170_),
    .X(_07314_));
 sky130_fd_sc_hd__buf_4 _12962_ (.A(_07165_),
    .X(_07315_));
 sky130_fd_sc_hd__a211o_1 _12963_ (.A1(_06606_),
    .A2(_06746_),
    .B1(_06790_),
    .C1(_06353_),
    .X(_07316_));
 sky130_fd_sc_hd__nand3_1 _12964_ (.A(_06353_),
    .B(_06407_),
    .C(_06607_),
    .Y(_07317_));
 sky130_fd_sc_hd__a21oi_1 _12965_ (.A1(_06407_),
    .A2(_06607_),
    .B1(_07165_),
    .Y(_07318_));
 sky130_fd_sc_hd__a31oi_1 _12966_ (.A1(_07315_),
    .A2(_07316_),
    .A3(_07317_),
    .B1(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_1 _12967_ (.A(net32),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(_06917_),
    .A1(_07040_),
    .S(_07164_),
    .X(_07321_));
 sky130_fd_sc_hd__clkbuf_4 _12969_ (.A(_07164_),
    .X(_07322_));
 sky130_fd_sc_hd__o221a_1 _12970_ (.A1(_06606_),
    .A2(_07062_),
    .B1(_07118_),
    .B2(_07161_),
    .C1(_06353_),
    .X(_07323_));
 sky130_fd_sc_hd__a311o_1 _12971_ (.A1(_07322_),
    .A2(_07201_),
    .A3(_07312_),
    .B1(_07323_),
    .C1(net31),
    .X(_07324_));
 sky130_fd_sc_hd__inv_2 _12972_ (.A(net32),
    .Y(_07325_));
 sky130_fd_sc_hd__clkbuf_4 _12973_ (.A(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__o211ai_4 _12974_ (.A1(_07315_),
    .A2(_07321_),
    .B1(_07324_),
    .C1(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__a21o_1 _12975_ (.A1(_06354_),
    .A2(_07167_),
    .B1(_07173_),
    .X(_07328_));
 sky130_fd_sc_hd__a31o_1 _12976_ (.A1(_07314_),
    .A2(_07320_),
    .A3(_07327_),
    .B1(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__or4_1 _12977_ (.A(_07165_),
    .B(_07164_),
    .C(_07170_),
    .D(_07325_),
    .X(_07330_));
 sky130_fd_sc_hd__buf_2 _12978_ (.A(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__o211a_2 _12979_ (.A1(_07182_),
    .A2(_07313_),
    .B1(_07329_),
    .C1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__xnor2_1 _12980_ (.A(\dsmod0.accu1[10] ),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__nor2_1 _12981_ (.A(_07180_),
    .B(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__mux4_1 _12982_ (.A0(\fifo0.fifo_store[76][9] ),
    .A1(\fifo0.fifo_store[77][9] ),
    .A2(\fifo0.fifo_store[78][9] ),
    .A3(\fifo0.fifo_store[79][9] ),
    .S0(_07097_),
    .S1(_06996_),
    .X(_07335_));
 sky130_fd_sc_hd__mux4_1 _12983_ (.A0(\fifo0.fifo_store[72][9] ),
    .A1(\fifo0.fifo_store[73][9] ),
    .A2(\fifo0.fifo_store[74][9] ),
    .A3(\fifo0.fifo_store[75][9] ),
    .S0(_06507_),
    .S1(_06975_),
    .X(_07336_));
 sky130_fd_sc_hd__or2_1 _12984_ (.A(_06474_),
    .B(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__o211a_1 _12985_ (.A1(_07071_),
    .A2(_07335_),
    .B1(_07337_),
    .C1(_07094_),
    .X(_07338_));
 sky130_fd_sc_hd__mux4_2 _12986_ (.A0(\fifo0.fifo_store[64][9] ),
    .A1(\fifo0.fifo_store[65][9] ),
    .A2(\fifo0.fifo_store[66][9] ),
    .A3(\fifo0.fifo_store[67][9] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_07339_));
 sky130_fd_sc_hd__or2b_1 _12987_ (.A(\fifo0.fifo_store[71][9] ),
    .B_N(_07067_),
    .X(_07340_));
 sky130_fd_sc_hd__o21a_1 _12988_ (.A1(_06416_),
    .A2(\fifo0.fifo_store[70][9] ),
    .B1(_06811_),
    .X(_07341_));
 sky130_fd_sc_hd__mux2_1 _12989_ (.A0(\fifo0.fifo_store[68][9] ),
    .A1(\fifo0.fifo_store[69][9] ),
    .S(_06956_),
    .X(_07342_));
 sky130_fd_sc_hd__a221o_1 _12990_ (.A1(_07340_),
    .A2(_07341_),
    .B1(_07342_),
    .B2(_07104_),
    .C1(_07132_),
    .X(_07343_));
 sky130_fd_sc_hd__o211a_1 _12991_ (.A1(_06442_),
    .A2(_07339_),
    .B1(_07343_),
    .C1(_06445_),
    .X(_07344_));
 sky130_fd_sc_hd__mux4_1 _12992_ (.A0(\fifo0.fifo_store[80][9] ),
    .A1(\fifo0.fifo_store[81][9] ),
    .A2(\fifo0.fifo_store[82][9] ),
    .A3(\fifo0.fifo_store[83][9] ),
    .S0(_06544_),
    .S1(_06695_),
    .X(_07345_));
 sky130_fd_sc_hd__mux4_1 _12993_ (.A0(\fifo0.fifo_store[84][9] ),
    .A1(\fifo0.fifo_store[85][9] ),
    .A2(\fifo0.fifo_store[86][9] ),
    .A3(\fifo0.fifo_store[87][9] ),
    .S0(_06544_),
    .S1(_06695_),
    .X(_07346_));
 sky130_fd_sc_hd__mux2_1 _12994_ (.A0(_07345_),
    .A1(_07346_),
    .S(_06730_),
    .X(_07347_));
 sky130_fd_sc_hd__mux4_1 _12995_ (.A0(\fifo0.fifo_store[88][9] ),
    .A1(\fifo0.fifo_store[89][9] ),
    .A2(\fifo0.fifo_store[90][9] ),
    .A3(\fifo0.fifo_store[91][9] ),
    .S0(_06697_),
    .S1(_07098_),
    .X(_07348_));
 sky130_fd_sc_hd__or2_1 _12996_ (.A(_06441_),
    .B(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__mux4_1 _12997_ (.A0(\fifo0.fifo_store[92][9] ),
    .A1(\fifo0.fifo_store[93][9] ),
    .A2(\fifo0.fifo_store[94][9] ),
    .A3(\fifo0.fifo_store[95][9] ),
    .S0(_06533_),
    .S1(_06592_),
    .X(_07350_));
 sky130_fd_sc_hd__o21a_1 _12998_ (.A1(_06517_),
    .A2(_07350_),
    .B1(_06462_),
    .X(_07351_));
 sky130_fd_sc_hd__a221o_1 _12999_ (.A1(_06445_),
    .A2(_07347_),
    .B1(_07349_),
    .B2(_07351_),
    .C1(_06539_),
    .X(_07352_));
 sky130_fd_sc_hd__o311a_1 _13000_ (.A1(_06409_),
    .A2(_07338_),
    .A3(_07344_),
    .B1(_07352_),
    .C1(_06498_),
    .X(_07353_));
 sky130_fd_sc_hd__buf_6 _13001_ (.A(_06539_),
    .X(_07354_));
 sky130_fd_sc_hd__buf_6 _13002_ (.A(_07132_),
    .X(_07355_));
 sky130_fd_sc_hd__mux4_1 _13003_ (.A0(\fifo0.fifo_store[124][9] ),
    .A1(\fifo0.fifo_store[125][9] ),
    .A2(\fifo0.fifo_store[126][9] ),
    .A3(\fifo0.fifo_store[127][9] ),
    .S0(_06435_),
    .S1(_06438_),
    .X(_07356_));
 sky130_fd_sc_hd__mux4_1 _13004_ (.A0(\fifo0.fifo_store[120][9] ),
    .A1(\fifo0.fifo_store[121][9] ),
    .A2(\fifo0.fifo_store[122][9] ),
    .A3(\fifo0.fifo_store[123][9] ),
    .S0(_06563_),
    .S1(_06561_),
    .X(_07357_));
 sky130_fd_sc_hd__or2_1 _13005_ (.A(_06797_),
    .B(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__o211a_1 _13006_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07358_),
    .C1(_06463_),
    .X(_07359_));
 sky130_fd_sc_hd__mux4_1 _13007_ (.A0(\fifo0.fifo_store[112][9] ),
    .A1(\fifo0.fifo_store[113][9] ),
    .A2(\fifo0.fifo_store[114][9] ),
    .A3(\fifo0.fifo_store[115][9] ),
    .S0(_06542_),
    .S1(_06454_),
    .X(_07360_));
 sky130_fd_sc_hd__or2b_1 _13008_ (.A(\fifo0.fifo_store[119][9] ),
    .B_N(_06545_),
    .X(_07361_));
 sky130_fd_sc_hd__o21a_1 _13009_ (.A1(_06545_),
    .A2(\fifo0.fifo_store[118][9] ),
    .B1(_06489_),
    .X(_07362_));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(\fifo0.fifo_store[116][9] ),
    .A1(\fifo0.fifo_store[117][9] ),
    .S(_07227_),
    .X(_07363_));
 sky130_fd_sc_hd__a221o_1 _13011_ (.A1(_07361_),
    .A2(_07362_),
    .B1(_07363_),
    .B2(_06516_),
    .C1(_06431_),
    .X(_07364_));
 sky130_fd_sc_hd__o211a_1 _13012_ (.A1(_06449_),
    .A2(_07360_),
    .B1(_07364_),
    .C1(_06468_),
    .X(_07365_));
 sky130_fd_sc_hd__mux4_2 _13013_ (.A0(\fifo0.fifo_store[96][9] ),
    .A1(\fifo0.fifo_store[97][9] ),
    .A2(\fifo0.fifo_store[98][9] ),
    .A3(\fifo0.fifo_store[99][9] ),
    .S0(_06434_),
    .S1(_07098_),
    .X(_07366_));
 sky130_fd_sc_hd__mux4_1 _13014_ (.A0(\fifo0.fifo_store[100][9] ),
    .A1(\fifo0.fifo_store[101][9] ),
    .A2(\fifo0.fifo_store[102][9] ),
    .A3(\fifo0.fifo_store[103][9] ),
    .S0(_06434_),
    .S1(_06561_),
    .X(_07367_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(_07366_),
    .A1(_07367_),
    .S(_06565_),
    .X(_07368_));
 sky130_fd_sc_hd__mux4_1 _13016_ (.A0(\fifo0.fifo_store[104][9] ),
    .A1(\fifo0.fifo_store[105][9] ),
    .A2(\fifo0.fifo_store[106][9] ),
    .A3(\fifo0.fifo_store[107][9] ),
    .S0(_06521_),
    .S1(_06523_),
    .X(_07369_));
 sky130_fd_sc_hd__or2_1 _13017_ (.A(_06519_),
    .B(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_6 _13018_ (.A(_06660_),
    .X(_07371_));
 sky130_fd_sc_hd__mux4_1 _13019_ (.A0(\fifo0.fifo_store[108][9] ),
    .A1(\fifo0.fifo_store[109][9] ),
    .A2(\fifo0.fifo_store[110][9] ),
    .A3(\fifo0.fifo_store[111][9] ),
    .S0(_07263_),
    .S1(_06481_),
    .X(_07372_));
 sky130_fd_sc_hd__o21a_1 _13020_ (.A1(_07371_),
    .A2(_07372_),
    .B1(_06571_),
    .X(_07373_));
 sky130_fd_sc_hd__a221o_1 _13021_ (.A1(_06552_),
    .A2(_07368_),
    .B1(_07370_),
    .B2(_07373_),
    .C1(_06589_),
    .X(_07374_));
 sky130_fd_sc_hd__o311a_1 _13022_ (.A1(_07354_),
    .A2(_07359_),
    .A3(_07365_),
    .B1(_06465_),
    .C1(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__nor3_4 _13023_ (.A(_06965_),
    .B(_07353_),
    .C(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__or2_1 _13024_ (.A(_06689_),
    .B(\fifo0.fifo_store[4][9] ),
    .X(_07377_));
 sky130_fd_sc_hd__o211a_1 _13025_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[5][9] ),
    .B1(_07377_),
    .C1(_06516_),
    .X(_07378_));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(\fifo0.fifo_store[6][9] ),
    .A1(\fifo0.fifo_store[7][9] ),
    .S(_06549_),
    .X(_07379_));
 sky130_fd_sc_hd__a21o_1 _13027_ (.A1(_07257_),
    .A2(_07379_),
    .B1(_06431_),
    .X(_07380_));
 sky130_fd_sc_hd__mux4_1 _13028_ (.A0(\fifo0.fifo_store[0][9] ),
    .A1(\fifo0.fifo_store[1][9] ),
    .A2(\fifo0.fifo_store[2][9] ),
    .A3(\fifo0.fifo_store[3][9] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_07381_));
 sky130_fd_sc_hd__o221ai_1 _13029_ (.A1(_07378_),
    .A2(_07380_),
    .B1(_07381_),
    .B2(_06442_),
    .C1(_06445_),
    .Y(_07382_));
 sky130_fd_sc_hd__mux4_1 _13030_ (.A0(\fifo0.fifo_store[12][9] ),
    .A1(\fifo0.fifo_store[13][9] ),
    .A2(\fifo0.fifo_store[14][9] ),
    .A3(\fifo0.fifo_store[15][9] ),
    .S0(_06452_),
    .S1(_06556_),
    .X(_07383_));
 sky130_fd_sc_hd__mux4_2 _13031_ (.A0(\fifo0.fifo_store[8][9] ),
    .A1(\fifo0.fifo_store[9][9] ),
    .A2(\fifo0.fifo_store[10][9] ),
    .A3(\fifo0.fifo_store[11][9] ),
    .S0(_06487_),
    .S1(_06489_),
    .X(_07384_));
 sky130_fd_sc_hd__o21a_1 _13032_ (.A1(_06485_),
    .A2(_07384_),
    .B1(_06491_),
    .X(_07385_));
 sky130_fd_sc_hd__o21ai_1 _13033_ (.A1(_07355_),
    .A2(_07383_),
    .B1(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__mux4_1 _13034_ (.A0(\fifo0.fifo_store[24][9] ),
    .A1(\fifo0.fifo_store[25][9] ),
    .A2(\fifo0.fifo_store[26][9] ),
    .A3(\fifo0.fifo_store[27][9] ),
    .S0(_06479_),
    .S1(_06811_),
    .X(_07387_));
 sky130_fd_sc_hd__nor2_1 _13035_ (.A(_06599_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__mux4_1 _13036_ (.A0(\fifo0.fifo_store[28][9] ),
    .A1(\fifo0.fifo_store[29][9] ),
    .A2(\fifo0.fifo_store[30][9] ),
    .A3(\fifo0.fifo_store[31][9] ),
    .S0(_06469_),
    .S1(_06471_),
    .X(_07389_));
 sky130_fd_sc_hd__o21ai_1 _13037_ (.A1(_06431_),
    .A2(_07389_),
    .B1(_06462_),
    .Y(_07390_));
 sky130_fd_sc_hd__clkbuf_16 _13038_ (.A(_06480_),
    .X(_07391_));
 sky130_fd_sc_hd__mux4_1 _13039_ (.A0(\fifo0.fifo_store[16][9] ),
    .A1(\fifo0.fifo_store[17][9] ),
    .A2(\fifo0.fifo_store[18][9] ),
    .A3(\fifo0.fifo_store[19][9] ),
    .S0(_07017_),
    .S1(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__nor2_1 _13040_ (.A(_06485_),
    .B(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__mux4_1 _13041_ (.A0(\fifo0.fifo_store[20][9] ),
    .A1(\fifo0.fifo_store[21][9] ),
    .A2(\fifo0.fifo_store[22][9] ),
    .A3(\fifo0.fifo_store[23][9] ),
    .S0(_06533_),
    .S1(_06592_),
    .X(_07394_));
 sky130_fd_sc_hd__o21ai_1 _13042_ (.A1(_06456_),
    .A2(_07394_),
    .B1(_06467_),
    .Y(_07395_));
 sky130_fd_sc_hd__o221a_1 _13043_ (.A1(_07388_),
    .A2(_07390_),
    .B1(_07393_),
    .B2(_07395_),
    .C1(_06408_),
    .X(_07396_));
 sky130_fd_sc_hd__a311o_1 _13044_ (.A1(_07085_),
    .A2(_07382_),
    .A3(_07386_),
    .B1(_06643_),
    .C1(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__or2_1 _13045_ (.A(_07001_),
    .B(\fifo0.fifo_store[52][9] ),
    .X(_07398_));
 sky130_fd_sc_hd__o211a_1 _13046_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[53][9] ),
    .B1(_07398_),
    .C1(_06425_),
    .X(_07399_));
 sky130_fd_sc_hd__mux2_1 _13047_ (.A0(\fifo0.fifo_store[54][9] ),
    .A1(\fifo0.fifo_store[55][9] ),
    .S(_07227_),
    .X(_07400_));
 sky130_fd_sc_hd__a21o_1 _13048_ (.A1(_06422_),
    .A2(_07400_),
    .B1(_06517_),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_1 _13049_ (.A0(\fifo0.fifo_store[48][9] ),
    .A1(\fifo0.fifo_store[49][9] ),
    .A2(\fifo0.fifo_store[50][9] ),
    .A3(\fifo0.fifo_store[51][9] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_07402_));
 sky130_fd_sc_hd__o221ai_4 _13050_ (.A1(_07399_),
    .A2(_07401_),
    .B1(_07402_),
    .B2(_06449_),
    .C1(_06552_),
    .Y(_07403_));
 sky130_fd_sc_hd__mux4_1 _13051_ (.A0(\fifo0.fifo_store[60][9] ),
    .A1(\fifo0.fifo_store[61][9] ),
    .A2(\fifo0.fifo_store[62][9] ),
    .A3(\fifo0.fifo_store[63][9] ),
    .S0(_06591_),
    .S1(_06592_),
    .X(_07404_));
 sky130_fd_sc_hd__nor2_1 _13052_ (.A(_06517_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__mux4_1 _13053_ (.A0(\fifo0.fifo_store[56][9] ),
    .A1(\fifo0.fifo_store[57][9] ),
    .A2(\fifo0.fifo_store[58][9] ),
    .A3(\fifo0.fifo_store[59][9] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_07406_));
 sky130_fd_sc_hd__nor2_1 _13054_ (.A(_06519_),
    .B(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__o31a_1 _13055_ (.A1(_06868_),
    .A2(_07405_),
    .A3(_07407_),
    .B1(_06641_),
    .X(_07408_));
 sky130_fd_sc_hd__mux4_1 _13056_ (.A0(\fifo0.fifo_store[36][9] ),
    .A1(\fifo0.fifo_store[37][9] ),
    .A2(\fifo0.fifo_store[38][9] ),
    .A3(\fifo0.fifo_store[39][9] ),
    .S0(_06499_),
    .S1(_06437_),
    .X(_07409_));
 sky130_fd_sc_hd__nor2_1 _13057_ (.A(_06517_),
    .B(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__mux4_1 _13058_ (.A0(\fifo0.fifo_store[32][9] ),
    .A1(\fifo0.fifo_store[33][9] ),
    .A2(\fifo0.fifo_store[34][9] ),
    .A3(\fifo0.fifo_store[35][9] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_07411_));
 sky130_fd_sc_hd__nor2_1 _13059_ (.A(_06448_),
    .B(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__mux4_1 _13060_ (.A0(\fifo0.fifo_store[40][9] ),
    .A1(\fifo0.fifo_store[41][9] ),
    .A2(\fifo0.fifo_store[42][9] ),
    .A3(\fifo0.fifo_store[43][9] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_07413_));
 sky130_fd_sc_hd__nor2_1 _13061_ (.A(_06624_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__mux4_1 _13062_ (.A0(\fifo0.fifo_store[44][9] ),
    .A1(\fifo0.fifo_store[45][9] ),
    .A2(\fifo0.fifo_store[46][9] ),
    .A3(\fifo0.fifo_store[47][9] ),
    .S0(_06810_),
    .S1(_06811_),
    .X(_07415_));
 sky130_fd_sc_hd__o21ai_1 _13063_ (.A1(_06477_),
    .A2(_07415_),
    .B1(_06491_),
    .Y(_07416_));
 sky130_fd_sc_hd__o32a_1 _13064_ (.A1(_06630_),
    .A2(_07410_),
    .A3(_07412_),
    .B1(_07414_),
    .B2(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__a221o_1 _13065_ (.A1(_07403_),
    .A2(_07408_),
    .B1(_07417_),
    .B2(_06679_),
    .C1(_06677_),
    .X(_07418_));
 sky130_fd_sc_hd__a31o_1 _13066_ (.A1(_06965_),
    .A2(_07397_),
    .A3(_07418_),
    .B1(_06918_),
    .X(_07419_));
 sky130_fd_sc_hd__a211o_1 _13067_ (.A1(_06378_),
    .A2(_06899_),
    .B1(_06368_),
    .C1(_06359_),
    .X(_07420_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(_06748_),
    .B(_06784_),
    .Y(_07421_));
 sky130_fd_sc_hd__nand2_1 _13069_ (.A(_06902_),
    .B(_06768_),
    .Y(_07422_));
 sky130_fd_sc_hd__a31o_1 _13070_ (.A1(_06378_),
    .A2(_07421_),
    .A3(_06779_),
    .B1(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__a21oi_1 _13071_ (.A1(_07420_),
    .A2(_07423_),
    .B1(_06370_),
    .Y(_07424_));
 sky130_fd_sc_hd__a31o_1 _13072_ (.A1(_06363_),
    .A2(_06751_),
    .A3(_06766_),
    .B1(_06373_),
    .X(_07425_));
 sky130_fd_sc_hd__or2b_1 _13073_ (.A(_07425_),
    .B_N(_06749_),
    .X(_07426_));
 sky130_fd_sc_hd__and3_1 _13074_ (.A(_06397_),
    .B(_06361_),
    .C(_06766_),
    .X(_07427_));
 sky130_fd_sc_hd__nor2_1 _13075_ (.A(_06912_),
    .B(_06361_),
    .Y(_07428_));
 sky130_fd_sc_hd__o21ai_1 _13076_ (.A1(_07427_),
    .A2(_07428_),
    .B1(_06359_),
    .Y(_07429_));
 sky130_fd_sc_hd__a31o_1 _13077_ (.A1(_06370_),
    .A2(_07426_),
    .A3(_07429_),
    .B1(_06769_),
    .X(_07430_));
 sky130_fd_sc_hd__o211a_1 _13078_ (.A1(_06391_),
    .A2(_06360_),
    .B1(_06766_),
    .C1(_06377_),
    .X(_07431_));
 sky130_fd_sc_hd__a211o_1 _13079_ (.A1(_06753_),
    .A2(_07431_),
    .B1(_06368_),
    .C1(_06902_),
    .X(_07432_));
 sky130_fd_sc_hd__a21o_1 _13080_ (.A1(_06922_),
    .A2(_06923_),
    .B1(_06401_),
    .X(_07433_));
 sky130_fd_sc_hd__a31o_1 _13081_ (.A1(_07421_),
    .A2(_06779_),
    .A3(_06893_),
    .B1(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__a311o_1 _13082_ (.A1(_06395_),
    .A2(_06398_),
    .A3(_06751_),
    .B1(_07184_),
    .C1(_06401_),
    .X(_07435_));
 sky130_fd_sc_hd__o21ba_2 _13083_ (.A1(_06390_),
    .A2(_06379_),
    .B1_N(_06376_),
    .X(_02165_));
 sky130_fd_sc_hd__a21o_1 _13084_ (.A1(_06399_),
    .A2(_02165_),
    .B1(_06373_),
    .X(_02166_));
 sky130_fd_sc_hd__and3_1 _13085_ (.A(_06397_),
    .B(_06384_),
    .C(_06784_),
    .X(_02167_));
 sky130_fd_sc_hd__o221a_1 _13086_ (.A1(_07427_),
    .A2(_07435_),
    .B1(_02166_),
    .B2(_02167_),
    .C1(_06369_),
    .X(_02168_));
 sky130_fd_sc_hd__a311o_1 _13087_ (.A1(_06405_),
    .A2(_07432_),
    .A3(_07434_),
    .B1(_02168_),
    .C1(_06919_),
    .X(_02169_));
 sky130_fd_sc_hd__o211ai_4 _13088_ (.A1(_07424_),
    .A2(_07430_),
    .B1(_06918_),
    .C1(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__o21ai_2 _13089_ (.A1(_07376_),
    .A2(_07419_),
    .B1(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__a211o_1 _13090_ (.A1(_06606_),
    .A2(_06746_),
    .B1(_06790_),
    .C1(_07163_),
    .X(_02172_));
 sky130_fd_sc_hd__a211o_1 _13091_ (.A1(_06841_),
    .A2(_06885_),
    .B1(_06916_),
    .C1(net30),
    .X(_02173_));
 sky130_fd_sc_hd__and2_1 _13092_ (.A(_02172_),
    .B(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__a2bb2o_1 _13093_ (.A1_N(_06991_),
    .A2_N(_07039_),
    .B1(_06918_),
    .B2(_06938_),
    .X(_02175_));
 sky130_fd_sc_hd__o22ai_1 _13094_ (.A1(_06611_),
    .A2(_07062_),
    .B1(_07118_),
    .B2(_07161_),
    .Y(_02176_));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(_02175_),
    .A1(_02176_),
    .S(_07164_),
    .X(_02177_));
 sky130_fd_sc_hd__o211a_1 _13096_ (.A1(_07376_),
    .A2(_07419_),
    .B1(_02170_),
    .C1(_07163_),
    .X(_02178_));
 sky130_fd_sc_hd__a31oi_2 _13097_ (.A1(_06353_),
    .A2(_07201_),
    .A3(_07312_),
    .B1(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__mux4_1 _13098_ (.A0(_07167_),
    .A1(_02174_),
    .A2(_02177_),
    .A3(_02179_),
    .S0(_07165_),
    .S1(_07325_),
    .X(_02180_));
 sky130_fd_sc_hd__a21o_1 _13099_ (.A1(_07314_),
    .A2(_02180_),
    .B1(_07328_),
    .X(_02181_));
 sky130_fd_sc_hd__o211a_1 _13100_ (.A1(_07182_),
    .A2(_02171_),
    .B1(_02181_),
    .C1(_07331_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_1 _13101_ (.A(\dsmod0.accu1[9] ),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__a21bo_1 _13102_ (.A1(_06693_),
    .A2(\fifo0.fifo_store[43][8] ),
    .B1_N(_06647_),
    .X(_02184_));
 sky130_fd_sc_hd__a21oi_1 _13103_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[42][8] ),
    .B1(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21o_1 _13104_ (.A1(_06549_),
    .A2(\fifo0.fifo_store[41][8] ),
    .B1(_06975_),
    .X(_02186_));
 sky130_fd_sc_hd__a21oi_1 _13105_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[40][8] ),
    .B1(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2b_1 _13106_ (.A(_06710_),
    .B_N(\fifo0.fifo_store[44][8] ),
    .X(_02188_));
 sky130_fd_sc_hd__a21oi_1 _13107_ (.A1(_06569_),
    .A2(\fifo0.fifo_store[45][8] ),
    .B1(_06984_),
    .Y(_02189_));
 sky130_fd_sc_hd__or2b_1 _13108_ (.A(_07008_),
    .B_N(\fifo0.fifo_store[46][8] ),
    .X(_02190_));
 sky130_fd_sc_hd__a21boi_1 _13109_ (.A1(_06487_),
    .A2(\fifo0.fifo_store[47][8] ),
    .B1_N(_06522_),
    .Y(_02191_));
 sky130_fd_sc_hd__a221o_1 _13110_ (.A1(_02188_),
    .A2(_02189_),
    .B1(_02190_),
    .B2(_02191_),
    .C1(_06430_),
    .X(_02192_));
 sky130_fd_sc_hd__o311a_1 _13111_ (.A1(_06474_),
    .A2(_02185_),
    .A3(_02187_),
    .B1(_02192_),
    .C1(_06462_),
    .X(_02193_));
 sky130_fd_sc_hd__and2_1 _13112_ (.A(_06617_),
    .B(\fifo0.fifo_store[35][8] ),
    .X(_02194_));
 sky130_fd_sc_hd__a211o_1 _13113_ (.A1(_06412_),
    .A2(\fifo0.fifo_store[34][8] ),
    .B1(_02194_),
    .C1(_06424_),
    .X(_02195_));
 sky130_fd_sc_hd__a21o_1 _13114_ (.A1(_06697_),
    .A2(\fifo0.fifo_store[33][8] ),
    .B1(_06510_),
    .X(_02196_));
 sky130_fd_sc_hd__a21o_1 _13115_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[32][8] ),
    .B1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__and2b_1 _13116_ (.A_N(_06617_),
    .B(\fifo0.fifo_store[36][8] ),
    .X(_02198_));
 sky130_fd_sc_hd__a21o_1 _13117_ (.A1(_07008_),
    .A2(\fifo0.fifo_store[37][8] ),
    .B1(_06522_),
    .X(_02199_));
 sky130_fd_sc_hd__and2b_1 _13118_ (.A_N(_06415_),
    .B(\fifo0.fifo_store[38][8] ),
    .X(_02200_));
 sky130_fd_sc_hd__a21bo_1 _13119_ (.A1(_06544_),
    .A2(\fifo0.fifo_store[39][8] ),
    .B1_N(_06470_),
    .X(_02201_));
 sky130_fd_sc_hd__o221a_1 _13120_ (.A1(_02198_),
    .A2(_02199_),
    .B1(_02200_),
    .B2(_02201_),
    .C1(_06447_),
    .X(_02202_));
 sky130_fd_sc_hd__a311o_1 _13121_ (.A1(_07132_),
    .A2(_02195_),
    .A3(_02197_),
    .B1(_06713_),
    .C1(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__or3b_1 _13122_ (.A(_06408_),
    .B(_02193_),
    .C_N(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__buf_6 _13123_ (.A(_06412_),
    .X(_02205_));
 sky130_fd_sc_hd__a21bo_1 _13124_ (.A1(_06870_),
    .A2(\fifo0.fifo_store[55][8] ),
    .B1_N(_06690_),
    .X(_02206_));
 sky130_fd_sc_hd__a21oi_1 _13125_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[54][8] ),
    .B1(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a21o_1 _13126_ (.A1(_06959_),
    .A2(\fifo0.fifo_store[53][8] ),
    .B1(_06561_),
    .X(_02208_));
 sky130_fd_sc_hd__a21oi_1 _13127_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[52][8] ),
    .B1(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__or2b_1 _13128_ (.A(_06507_),
    .B_N(\fifo0.fifo_store[50][8] ),
    .X(_02210_));
 sky130_fd_sc_hd__a21boi_1 _13129_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[51][8] ),
    .B1_N(_06488_),
    .Y(_02211_));
 sky130_fd_sc_hd__or2b_1 _13130_ (.A(_06645_),
    .B_N(\fifo0.fifo_store[48][8] ),
    .X(_02212_));
 sky130_fd_sc_hd__a21oi_1 _13131_ (.A1(_06549_),
    .A2(\fifo0.fifo_store[49][8] ),
    .B1(_06975_),
    .Y(_02213_));
 sky130_fd_sc_hd__a221o_1 _13132_ (.A1(_02210_),
    .A2(_02211_),
    .B1(_02212_),
    .B2(_02213_),
    .C1(_06447_),
    .X(_02214_));
 sky130_fd_sc_hd__o311a_1 _13133_ (.A1(_07132_),
    .A2(_02207_),
    .A3(_02209_),
    .B1(_06467_),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__a21bo_1 _13134_ (.A1(_06514_),
    .A2(\fifo0.fifo_store[59][8] ),
    .B1_N(_06711_),
    .X(_02216_));
 sky130_fd_sc_hd__a21oi_1 _13135_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[58][8] ),
    .B1(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__a21o_1 _13136_ (.A1(_06689_),
    .A2(\fifo0.fifo_store[57][8] ),
    .B1(_06471_),
    .X(_02218_));
 sky130_fd_sc_hd__a21oi_1 _13137_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[56][8] ),
    .B1(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__or2b_1 _13138_ (.A(_06527_),
    .B_N(\fifo0.fifo_store[60][8] ),
    .X(_02220_));
 sky130_fd_sc_hd__a21oi_1 _13139_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[61][8] ),
    .B1(_06975_),
    .Y(_02221_));
 sky130_fd_sc_hd__or2b_1 _13140_ (.A(_06645_),
    .B_N(\fifo0.fifo_store[62][8] ),
    .X(_02222_));
 sky130_fd_sc_hd__a21boi_1 _13141_ (.A1(_06549_),
    .A2(\fifo0.fifo_store[63][8] ),
    .B1_N(_06578_),
    .Y(_02223_));
 sky130_fd_sc_hd__a221o_1 _13142_ (.A1(_02220_),
    .A2(_02221_),
    .B1(_02222_),
    .B2(_02223_),
    .C1(_06476_),
    .X(_02224_));
 sky130_fd_sc_hd__o311a_1 _13143_ (.A1(_06448_),
    .A2(_02217_),
    .A3(_02219_),
    .B1(_02224_),
    .C1(_07219_),
    .X(_02225_));
 sky130_fd_sc_hd__o31a_2 _13144_ (.A1(_06539_),
    .A2(_02215_),
    .A3(_02225_),
    .B1(_00005_),
    .X(_02226_));
 sky130_fd_sc_hd__and2_1 _13145_ (.A(_06870_),
    .B(\fifo0.fifo_store[31][8] ),
    .X(_02227_));
 sky130_fd_sc_hd__a211o_1 _13146_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[30][8] ),
    .B1(_02227_),
    .C1(_07104_),
    .X(_02228_));
 sky130_fd_sc_hd__a21o_1 _13147_ (.A1(_06545_),
    .A2(\fifo0.fifo_store[29][8] ),
    .B1(_06811_),
    .X(_02229_));
 sky130_fd_sc_hd__a21o_1 _13148_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[28][8] ),
    .B1(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__and3_1 _13149_ (.A(_06688_),
    .B(_02228_),
    .C(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__and2_1 _13150_ (.A(_07022_),
    .B(\fifo0.fifo_store[27][8] ),
    .X(_02232_));
 sky130_fd_sc_hd__a211o_1 _13151_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[26][8] ),
    .B1(_02232_),
    .C1(_07104_),
    .X(_02233_));
 sky130_fd_sc_hd__buf_6 _13152_ (.A(_06412_),
    .X(_02234_));
 sky130_fd_sc_hd__a21o_1 _13153_ (.A1(_07097_),
    .A2(\fifo0.fifo_store[25][8] ),
    .B1(_06579_),
    .X(_02235_));
 sky130_fd_sc_hd__a21o_1 _13154_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[24][8] ),
    .B1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__a31o_1 _13155_ (.A1(_07071_),
    .A2(_02233_),
    .A3(_02236_),
    .B1(_07107_),
    .X(_02237_));
 sky130_fd_sc_hd__and2_1 _13156_ (.A(_07227_),
    .B(\fifo0.fifo_store[19][8] ),
    .X(_02238_));
 sky130_fd_sc_hd__a211o_1 _13157_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[18][8] ),
    .B1(_02238_),
    .C1(_07104_),
    .X(_02239_));
 sky130_fd_sc_hd__a21o_1 _13158_ (.A1(_06576_),
    .A2(\fifo0.fifo_store[17][8] ),
    .B1(_07391_),
    .X(_02240_));
 sky130_fd_sc_hd__a21o_1 _13159_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[16][8] ),
    .B1(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__and2b_1 _13160_ (.A_N(_06514_),
    .B(\fifo0.fifo_store[20][8] ),
    .X(_02242_));
 sky130_fd_sc_hd__a21o_1 _13161_ (.A1(_06689_),
    .A2(\fifo0.fifo_store[21][8] ),
    .B1(_06437_),
    .X(_02243_));
 sky130_fd_sc_hd__and2b_1 _13162_ (.A_N(_06959_),
    .B(\fifo0.fifo_store[22][8] ),
    .X(_02244_));
 sky130_fd_sc_hd__a21bo_1 _13163_ (.A1(_06416_),
    .A2(\fifo0.fifo_store[23][8] ),
    .B1_N(_07111_),
    .X(_02245_));
 sky130_fd_sc_hd__o221a_1 _13164_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02244_),
    .B2(_02245_),
    .C1(_06797_),
    .X(_02246_));
 sky130_fd_sc_hd__a311o_1 _13165_ (.A1(_07071_),
    .A2(_02239_),
    .A3(_02241_),
    .B1(_06686_),
    .C1(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__o211ai_1 _13166_ (.A1(_02231_),
    .A2(_02237_),
    .B1(_06409_),
    .C1(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__a21bo_1 _13167_ (.A1(_06427_),
    .A2(\fifo0.fifo_store[11][8] ),
    .B1_N(_06984_),
    .X(_02249_));
 sky130_fd_sc_hd__a21oi_2 _13168_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[10][8] ),
    .B1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21o_1 _13169_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[9][8] ),
    .B1(_07098_),
    .X(_02251_));
 sky130_fd_sc_hd__a21oi_1 _13170_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[8][8] ),
    .B1(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__or2b_1 _13171_ (.A(_06507_),
    .B_N(\fifo0.fifo_store[12][8] ),
    .X(_02253_));
 sky130_fd_sc_hd__a21oi_1 _13172_ (.A1(_06956_),
    .A2(\fifo0.fifo_store[13][8] ),
    .B1(_06695_),
    .Y(_02254_));
 sky130_fd_sc_hd__or2b_1 _13173_ (.A(_06507_),
    .B_N(\fifo0.fifo_store[14][8] ),
    .X(_02255_));
 sky130_fd_sc_hd__a21boi_1 _13174_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[15][8] ),
    .B1_N(_06488_),
    .Y(_02256_));
 sky130_fd_sc_hd__a221o_1 _13175_ (.A1(_02253_),
    .A2(_02254_),
    .B1(_02255_),
    .B2(_02256_),
    .C1(_06476_),
    .X(_02257_));
 sky130_fd_sc_hd__o311a_1 _13176_ (.A1(_06441_),
    .A2(_02250_),
    .A3(_02252_),
    .B1(_02257_),
    .C1(_06491_),
    .X(_02258_));
 sky130_fd_sc_hd__a21bo_1 _13177_ (.A1(_06959_),
    .A2(\fifo0.fifo_store[3][8] ),
    .B1_N(_06725_),
    .X(_02259_));
 sky130_fd_sc_hd__a21oi_1 _13178_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[2][8] ),
    .B1(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21o_1 _13179_ (.A1(_06689_),
    .A2(\fifo0.fifo_store[1][8] ),
    .B1(_06592_),
    .X(_02261_));
 sky130_fd_sc_hd__a21oi_1 _13180_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[0][8] ),
    .B1(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__or2b_1 _13181_ (.A(_06697_),
    .B_N(\fifo0.fifo_store[4][8] ),
    .X(_02263_));
 sky130_fd_sc_hd__a21oi_1 _13182_ (.A1(_06514_),
    .A2(\fifo0.fifo_store[5][8] ),
    .B1(_06561_),
    .Y(_02264_));
 sky130_fd_sc_hd__buf_8 _13183_ (.A(_06414_),
    .X(_02265_));
 sky130_fd_sc_hd__or2b_1 _13184_ (.A(_02265_),
    .B_N(\fifo0.fifo_store[6][8] ),
    .X(_02266_));
 sky130_fd_sc_hd__a21boi_1 _13185_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[7][8] ),
    .B1_N(_06614_),
    .Y(_02267_));
 sky130_fd_sc_hd__a221o_1 _13186_ (.A1(_02263_),
    .A2(_02264_),
    .B1(_02266_),
    .B2(_02267_),
    .C1(_06660_),
    .X(_02268_));
 sky130_fd_sc_hd__o311a_1 _13187_ (.A1(_06448_),
    .A2(_02260_),
    .A3(_02262_),
    .B1(_06621_),
    .C1(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__o31a_1 _13188_ (.A1(_06589_),
    .A2(_02258_),
    .A3(_02269_),
    .B1(_06497_),
    .X(_02270_));
 sky130_fd_sc_hd__a221o_4 _13189_ (.A1(_02204_),
    .A2(_02226_),
    .B1(_02248_),
    .B2(_02270_),
    .C1(_00006_),
    .X(_02271_));
 sky130_fd_sc_hd__and2_1 _13190_ (.A(_06569_),
    .B(\fifo0.fifo_store[107][8] ),
    .X(_02272_));
 sky130_fd_sc_hd__a211o_1 _13191_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[106][8] ),
    .B1(_02272_),
    .C1(_06728_),
    .X(_02273_));
 sky130_fd_sc_hd__a21o_1 _13192_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[105][8] ),
    .B1(_07098_),
    .X(_02274_));
 sky130_fd_sc_hd__a21o_1 _13193_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[104][8] ),
    .B1(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__and2b_1 _13194_ (.A_N(_07263_),
    .B(\fifo0.fifo_store[110][8] ),
    .X(_02276_));
 sky130_fd_sc_hd__a21bo_1 _13195_ (.A1(_06658_),
    .A2(\fifo0.fifo_store[111][8] ),
    .B1_N(_06731_),
    .X(_02277_));
 sky130_fd_sc_hd__and2b_1 _13196_ (.A_N(_06487_),
    .B(\fifo0.fifo_store[108][8] ),
    .X(_02278_));
 sky130_fd_sc_hd__a21o_1 _13197_ (.A1(_06549_),
    .A2(\fifo0.fifo_store[109][8] ),
    .B1(_06975_),
    .X(_02279_));
 sky130_fd_sc_hd__o221a_1 _13198_ (.A1(_02276_),
    .A2(_02277_),
    .B1(_02278_),
    .B2(_02279_),
    .C1(_06531_),
    .X(_02280_));
 sky130_fd_sc_hd__a311o_1 _13199_ (.A1(_06945_),
    .A2(_02273_),
    .A3(_02275_),
    .B1(_06735_),
    .C1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__and2_1 _13200_ (.A(_06479_),
    .B(\fifo0.fifo_store[99][8] ),
    .X(_02282_));
 sky130_fd_sc_hd__a211o_1 _13201_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[98][8] ),
    .B1(_02282_),
    .C1(_06728_),
    .X(_02283_));
 sky130_fd_sc_hd__a21o_1 _13202_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[97][8] ),
    .B1(_07098_),
    .X(_02284_));
 sky130_fd_sc_hd__a21o_1 _13203_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[96][8] ),
    .B1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__and2b_1 _13204_ (.A_N(_07263_),
    .B(\fifo0.fifo_store[100][8] ),
    .X(_02286_));
 sky130_fd_sc_hd__a21o_1 _13205_ (.A1(_06956_),
    .A2(\fifo0.fifo_store[101][8] ),
    .B1(_06695_),
    .X(_02287_));
 sky130_fd_sc_hd__and2b_1 _13206_ (.A_N(_06487_),
    .B(\fifo0.fifo_store[102][8] ),
    .X(_02288_));
 sky130_fd_sc_hd__a21bo_1 _13207_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[103][8] ),
    .B1_N(_06690_),
    .X(_02289_));
 sky130_fd_sc_hd__o221a_1 _13208_ (.A1(_02286_),
    .A2(_02287_),
    .B1(_02288_),
    .B2(_02289_),
    .C1(_06730_),
    .X(_02290_));
 sky130_fd_sc_hd__a311o_1 _13209_ (.A1(_06681_),
    .A2(_02283_),
    .A3(_02285_),
    .B1(_06664_),
    .C1(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__and3_1 _13210_ (.A(_07085_),
    .B(_02281_),
    .C(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__and2_1 _13211_ (.A(_06693_),
    .B(\fifo0.fifo_store[115][8] ),
    .X(_02293_));
 sky130_fd_sc_hd__a211o_1 _13212_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[114][8] ),
    .B1(_02293_),
    .C1(_06699_),
    .X(_02294_));
 sky130_fd_sc_hd__a21o_1 _13213_ (.A1(_07001_),
    .A2(\fifo0.fifo_store[113][8] ),
    .B1(_06458_),
    .X(_02295_));
 sky130_fd_sc_hd__a21o_1 _13214_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[112][8] ),
    .B1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__and2b_1 _13215_ (.A_N(_06848_),
    .B(\fifo0.fifo_store[116][8] ),
    .X(_02297_));
 sky130_fd_sc_hd__a21o_1 _13216_ (.A1(_07227_),
    .A2(\fifo0.fifo_store[117][8] ),
    .B1(_07111_),
    .X(_02298_));
 sky130_fd_sc_hd__and2b_1 _13217_ (.A_N(_06801_),
    .B(\fifo0.fifo_store[118][8] ),
    .X(_02299_));
 sky130_fd_sc_hd__a21bo_1 _13218_ (.A1(_06514_),
    .A2(\fifo0.fifo_store[119][8] ),
    .B1_N(_06711_),
    .X(_02300_));
 sky130_fd_sc_hd__o221a_1 _13219_ (.A1(_02297_),
    .A2(_02298_),
    .B1(_02299_),
    .B2(_02300_),
    .C1(_06565_),
    .X(_02301_));
 sky130_fd_sc_hd__a311o_1 _13220_ (.A1(_06945_),
    .A2(_02294_),
    .A3(_02296_),
    .B1(_06664_),
    .C1(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__a21o_1 _13221_ (.A1(_06416_),
    .A2(\fifo0.fifo_store[125][8] ),
    .B1(_06453_),
    .X(_02303_));
 sky130_fd_sc_hd__a21o_1 _13222_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[124][8] ),
    .B1(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(_06625_),
    .B(\fifo0.fifo_store[127][8] ),
    .X(_02305_));
 sky130_fd_sc_hd__a211o_1 _13224_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[126][8] ),
    .B1(_02305_),
    .C1(_06699_),
    .X(_02306_));
 sky130_fd_sc_hd__and2b_1 _13225_ (.A_N(_06848_),
    .B(\fifo0.fifo_store[122][8] ),
    .X(_02307_));
 sky130_fd_sc_hd__a21bo_1 _13226_ (.A1(_06427_),
    .A2(\fifo0.fifo_store[123][8] ),
    .B1_N(_06984_),
    .X(_02308_));
 sky130_fd_sc_hd__and2b_1 _13227_ (.A_N(_06956_),
    .B(\fifo0.fifo_store[120][8] ),
    .X(_02309_));
 sky130_fd_sc_hd__a21o_1 _13228_ (.A1(_06959_),
    .A2(\fifo0.fifo_store[121][8] ),
    .B1(_06561_),
    .X(_02310_));
 sky130_fd_sc_hd__o221a_1 _13229_ (.A1(_02307_),
    .A2(_02308_),
    .B1(_02309_),
    .B2(_02310_),
    .C1(_06721_),
    .X(_02311_));
 sky130_fd_sc_hd__a311o_1 _13230_ (.A1(_06688_),
    .A2(_02304_),
    .A3(_02306_),
    .B1(_06701_),
    .C1(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__a31o_1 _13231_ (.A1(_06966_),
    .A2(_02302_),
    .A3(_02312_),
    .B1(_06498_),
    .X(_02313_));
 sky130_fd_sc_hd__a21o_1 _13232_ (.A1(_06689_),
    .A2(\fifo0.fifo_store[85][8] ),
    .B1(_06437_),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _13233_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[84][8] ),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__and2_1 _13234_ (.A(_07017_),
    .B(\fifo0.fifo_store[87][8] ),
    .X(_02316_));
 sky130_fd_sc_hd__a211o_1 _13235_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[86][8] ),
    .B1(_02316_),
    .C1(_06699_),
    .X(_02317_));
 sky130_fd_sc_hd__and2b_1 _13236_ (.A_N(_06487_),
    .B(\fifo0.fifo_store[80][8] ),
    .X(_02318_));
 sky130_fd_sc_hd__a21o_1 _13237_ (.A1(_06870_),
    .A2(\fifo0.fifo_store[81][8] ),
    .B1(_07072_),
    .X(_02319_));
 sky130_fd_sc_hd__and2b_1 _13238_ (.A_N(_06848_),
    .B(\fifo0.fifo_store[82][8] ),
    .X(_02320_));
 sky130_fd_sc_hd__a21bo_1 _13239_ (.A1(_06427_),
    .A2(\fifo0.fifo_store[83][8] ),
    .B1_N(_06984_),
    .X(_02321_));
 sky130_fd_sc_hd__o221a_1 _13240_ (.A1(_02318_),
    .A2(_02319_),
    .B1(_02320_),
    .B2(_02321_),
    .C1(_06721_),
    .X(_02322_));
 sky130_fd_sc_hd__a311o_1 _13241_ (.A1(_06688_),
    .A2(_02315_),
    .A3(_02317_),
    .B1(_06664_),
    .C1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__and2_1 _13242_ (.A(_07017_),
    .B(\fifo0.fifo_store[91][8] ),
    .X(_02324_));
 sky130_fd_sc_hd__a211o_1 _13243_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[90][8] ),
    .B1(_02324_),
    .C1(_06699_),
    .X(_02325_));
 sky130_fd_sc_hd__a21o_1 _13244_ (.A1(_06689_),
    .A2(\fifo0.fifo_store[89][8] ),
    .B1(_06471_),
    .X(_02326_));
 sky130_fd_sc_hd__a21o_1 _13245_ (.A1(_07226_),
    .A2(\fifo0.fifo_store[88][8] ),
    .B1(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__and2b_1 _13246_ (.A_N(_06487_),
    .B(\fifo0.fifo_store[94][8] ),
    .X(_02328_));
 sky130_fd_sc_hd__a21bo_1 _13247_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[95][8] ),
    .B1_N(_06690_),
    .X(_02329_));
 sky130_fd_sc_hd__and2b_1 _13248_ (.A_N(_06848_),
    .B(\fifo0.fifo_store[92][8] ),
    .X(_02330_));
 sky130_fd_sc_hd__a21o_1 _13249_ (.A1(_07227_),
    .A2(\fifo0.fifo_store[93][8] ),
    .B1(_06528_),
    .X(_02331_));
 sky130_fd_sc_hd__o221a_1 _13250_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02330_),
    .B2(_02331_),
    .C1(_06531_),
    .X(_02332_));
 sky130_fd_sc_hd__a311o_1 _13251_ (.A1(_06945_),
    .A2(_02325_),
    .A3(_02327_),
    .B1(_06735_),
    .C1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__and3_1 _13252_ (.A(_06966_),
    .B(_02323_),
    .C(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__a21o_1 _13253_ (.A1(_07067_),
    .A2(\fifo0.fifo_store[77][8] ),
    .B1(_06555_),
    .X(_02335_));
 sky130_fd_sc_hd__a21o_1 _13254_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[76][8] ),
    .B1(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__and2_1 _13255_ (.A(_06956_),
    .B(\fifo0.fifo_store[79][8] ),
    .X(_02337_));
 sky130_fd_sc_hd__a211o_1 _13256_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[78][8] ),
    .B1(_02337_),
    .C1(_06699_),
    .X(_02338_));
 sky130_fd_sc_hd__and2b_1 _13257_ (.A_N(_06870_),
    .B(\fifo0.fifo_store[72][8] ),
    .X(_02339_));
 sky130_fd_sc_hd__a21o_1 _13258_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[73][8] ),
    .B1(_07098_),
    .X(_02340_));
 sky130_fd_sc_hd__and2b_1 _13259_ (.A_N(_06427_),
    .B(\fifo0.fifo_store[74][8] ),
    .X(_02341_));
 sky130_fd_sc_hd__a21bo_1 _13260_ (.A1(_06946_),
    .A2(\fifo0.fifo_store[75][8] ),
    .B1_N(_07072_),
    .X(_02342_));
 sky130_fd_sc_hd__o221a_1 _13261_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02341_),
    .B2(_02342_),
    .C1(_06709_),
    .X(_02343_));
 sky130_fd_sc_hd__a311o_1 _13262_ (.A1(_07066_),
    .A2(_02336_),
    .A3(_02338_),
    .B1(_06701_),
    .C1(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__and2_1 _13263_ (.A(_06956_),
    .B(\fifo0.fifo_store[67][8] ),
    .X(_02345_));
 sky130_fd_sc_hd__a211o_1 _13264_ (.A1(_07119_),
    .A2(\fifo0.fifo_store[66][8] ),
    .B1(_02345_),
    .C1(_06699_),
    .X(_02346_));
 sky130_fd_sc_hd__a21o_1 _13265_ (.A1(_07067_),
    .A2(\fifo0.fifo_store[65][8] ),
    .B1(_06523_),
    .X(_02347_));
 sky130_fd_sc_hd__a21o_1 _13266_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[64][8] ),
    .B1(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__and2b_1 _13267_ (.A_N(_06870_),
    .B(\fifo0.fifo_store[68][8] ),
    .X(_02349_));
 sky130_fd_sc_hd__a21o_1 _13268_ (.A1(_07022_),
    .A2(\fifo0.fifo_store[69][8] ),
    .B1(_07098_),
    .X(_02350_));
 sky130_fd_sc_hd__and2b_1 _13269_ (.A_N(_06427_),
    .B(\fifo0.fifo_store[70][8] ),
    .X(_02351_));
 sky130_fd_sc_hd__a21bo_1 _13270_ (.A1(_06946_),
    .A2(\fifo0.fifo_store[71][8] ),
    .B1_N(_07072_),
    .X(_02352_));
 sky130_fd_sc_hd__o221a_1 _13271_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_02351_),
    .B2(_02352_),
    .C1(_06474_),
    .X(_02353_));
 sky130_fd_sc_hd__a311o_1 _13272_ (.A1(_06945_),
    .A2(_02346_),
    .A3(_02348_),
    .B1(_06686_),
    .C1(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__a31o_1 _13273_ (.A1(_07085_),
    .A2(_02344_),
    .A3(_02354_),
    .B1(_06643_),
    .X(_02355_));
 sky130_fd_sc_hd__o221ai_4 _13274_ (.A1(_02292_),
    .A2(_02313_),
    .B1(_02334_),
    .B2(_02355_),
    .C1(_06992_),
    .Y(_02356_));
 sky130_fd_sc_hd__o221a_1 _13275_ (.A1(_06397_),
    .A2(_06386_),
    .B1(_06759_),
    .B2(_06748_),
    .C1(_06401_),
    .X(_02357_));
 sky130_fd_sc_hd__nor2_1 _13276_ (.A(_06377_),
    .B(_06399_),
    .Y(_02358_));
 sky130_fd_sc_hd__o311a_1 _13277_ (.A1(_06382_),
    .A2(_06774_),
    .A3(_02358_),
    .B1(_06768_),
    .C1(_06358_),
    .X(_02359_));
 sky130_fd_sc_hd__a311o_1 _13278_ (.A1(_06761_),
    .A2(_06775_),
    .A3(_02357_),
    .B1(_02359_),
    .C1(_06369_),
    .X(_02360_));
 sky130_fd_sc_hd__o31ai_1 _13279_ (.A1(_06359_),
    .A2(_06911_),
    .A3(_07052_),
    .B1(_06370_),
    .Y(_02361_));
 sky130_fd_sc_hd__a32o_1 _13280_ (.A1(_06378_),
    .A2(_06751_),
    .A3(_06766_),
    .B1(_06891_),
    .B2(_06784_),
    .X(_02362_));
 sky130_fd_sc_hd__a221o_1 _13281_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02362_),
    .B2(_06910_),
    .C1(_06919_),
    .X(_02363_));
 sky130_fd_sc_hd__a221o_1 _13282_ (.A1(_06924_),
    .A2(_06922_),
    .B1(_07058_),
    .B2(_07057_),
    .C1(_06374_),
    .X(_02364_));
 sky130_fd_sc_hd__nand3_1 _13283_ (.A(_06399_),
    .B(_02165_),
    .C(_06753_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21oi_1 _13284_ (.A1(_06772_),
    .A2(_02365_),
    .B1(_06902_),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _13285_ (.A(_06910_),
    .Y(_02367_));
 sky130_fd_sc_hd__o32a_1 _13286_ (.A1(_06370_),
    .A2(_02359_),
    .A3(_02366_),
    .B1(_02362_),
    .B2(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__a31oi_2 _13287_ (.A1(_06919_),
    .A2(_02364_),
    .A3(_02368_),
    .B1(_06357_),
    .Y(_02369_));
 sky130_fd_sc_hd__a32oi_4 _13288_ (.A1(_06606_),
    .A2(_02271_),
    .A3(_02356_),
    .B1(_02363_),
    .B2(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__a21o_1 _13289_ (.A1(_06841_),
    .A2(_06885_),
    .B1(_06916_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _13290_ (.A0(_02371_),
    .A1(_02175_),
    .S(_07163_),
    .X(_02372_));
 sky130_fd_sc_hd__and2_1 _13291_ (.A(_07316_),
    .B(_07317_),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(_02171_),
    .A1(_02370_),
    .S(_07163_),
    .X(_02374_));
 sky130_fd_sc_hd__a31oi_1 _13293_ (.A1(_07164_),
    .A2(_07201_),
    .A3(_07312_),
    .B1(_07323_),
    .Y(_02375_));
 sky130_fd_sc_hd__mux4_1 _13294_ (.A0(_02372_),
    .A1(_02373_),
    .A2(_02374_),
    .A3(_02375_),
    .S0(net31),
    .S1(_07326_),
    .X(_02376_));
 sky130_fd_sc_hd__a21o_1 _13295_ (.A1(_07314_),
    .A2(_02376_),
    .B1(_07328_),
    .X(_02377_));
 sky130_fd_sc_hd__o211a_1 _13296_ (.A1(_07182_),
    .A2(_02370_),
    .B1(_02377_),
    .C1(_07331_),
    .X(_02378_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(\dsmod0.accu1[8] ),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__nor2_1 _13298_ (.A(\dsmod0.accu1[9] ),
    .B(_02182_),
    .Y(_02380_));
 sky130_fd_sc_hd__a21oi_1 _13299_ (.A1(_02183_),
    .A2(_02379_),
    .B1(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__inv_2 _13300_ (.A(\dsmod0.accu1[5] ),
    .Y(_02382_));
 sky130_fd_sc_hd__buf_2 _13301_ (.A(_07331_),
    .X(_02383_));
 sky130_fd_sc_hd__a31o_1 _13302_ (.A1(_07315_),
    .A2(_02172_),
    .A3(_02173_),
    .B1(_07318_),
    .X(_02384_));
 sky130_fd_sc_hd__a21bo_1 _13303_ (.A1(_07326_),
    .A2(_02384_),
    .B1_N(_07168_),
    .X(_02385_));
 sky130_fd_sc_hd__o21ai_1 _13304_ (.A1(_06762_),
    .A2(_06899_),
    .B1(_07195_),
    .Y(_02386_));
 sky130_fd_sc_hd__a2111o_1 _13305_ (.A1(_06397_),
    .A2(_06382_),
    .B1(_02358_),
    .C1(_06380_),
    .D1(_06401_),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _13306_ (.A(_06369_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__a21oi_1 _13307_ (.A1(_06402_),
    .A2(_02386_),
    .B1(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand3_1 _13308_ (.A(_06373_),
    .B(_06399_),
    .C(_02165_),
    .Y(_02390_));
 sky130_fd_sc_hd__o31a_1 _13309_ (.A1(_06401_),
    .A2(_06393_),
    .A3(_06920_),
    .B1(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__o311a_1 _13310_ (.A1(_06902_),
    .A2(_06903_),
    .A3(_06762_),
    .B1(_02391_),
    .C1(_06404_),
    .X(_02392_));
 sky130_fd_sc_hd__o21a_1 _13311_ (.A1(_02389_),
    .A2(_02392_),
    .B1(_06769_),
    .X(_02393_));
 sky130_fd_sc_hd__a211o_1 _13312_ (.A1(_06378_),
    .A2(_06384_),
    .B1(_06762_),
    .C1(_06358_),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_1 _13313_ (.A(_02391_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(_06396_),
    .B(_06899_),
    .Y(_02396_));
 sky130_fd_sc_hd__o21a_1 _13315_ (.A1(_06913_),
    .A2(_02396_),
    .B1(_06402_),
    .X(_02397_));
 sky130_fd_sc_hd__o221a_1 _13316_ (.A1(_06370_),
    .A2(_02395_),
    .B1(_02397_),
    .B2(_02388_),
    .C1(_06919_),
    .X(_02398_));
 sky130_fd_sc_hd__buf_4 _13317_ (.A(_06412_),
    .X(_02399_));
 sky130_fd_sc_hd__and2_1 _13318_ (.A(_06586_),
    .B(\fifo0.fifo_store[43][7] ),
    .X(_02400_));
 sky130_fd_sc_hd__a211o_1 _13319_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[42][7] ),
    .B1(_02400_),
    .C1(_06650_),
    .X(_02401_));
 sky130_fd_sc_hd__a21o_1 _13320_ (.A1(_06658_),
    .A2(\fifo0.fifo_store[41][7] ),
    .B1(_06725_),
    .X(_02402_));
 sky130_fd_sc_hd__a21o_1 _13321_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[40][7] ),
    .B1(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__and3_1 _13322_ (.A(_07371_),
    .B(_02401_),
    .C(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__a21o_1 _13323_ (.A1(_06870_),
    .A2(\fifo0.fifo_store[45][7] ),
    .B1(_06975_),
    .X(_02405_));
 sky130_fd_sc_hd__a21o_1 _13324_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[44][7] ),
    .B1(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__clkbuf_8 _13325_ (.A(_06412_),
    .X(_02407_));
 sky130_fd_sc_hd__and2_1 _13326_ (.A(_06499_),
    .B(\fifo0.fifo_store[47][7] ),
    .X(_02408_));
 sky130_fd_sc_hd__a211o_1 _13327_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[46][7] ),
    .B1(_02408_),
    .C1(_06829_),
    .X(_02409_));
 sky130_fd_sc_hd__a31o_1 _13328_ (.A1(_06656_),
    .A2(_02406_),
    .A3(_02409_),
    .B1(_06621_),
    .X(_02410_));
 sky130_fd_sc_hd__a21o_1 _13329_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[37][7] ),
    .B1(_07072_),
    .X(_02411_));
 sky130_fd_sc_hd__a21o_1 _13330_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[36][7] ),
    .B1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__and2_1 _13331_ (.A(_02265_),
    .B(\fifo0.fifo_store[39][7] ),
    .X(_02413_));
 sky130_fd_sc_hd__a211o_1 _13332_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[38][7] ),
    .B1(_02413_),
    .C1(_06829_),
    .X(_02414_));
 sky130_fd_sc_hd__and3_1 _13333_ (.A(_06624_),
    .B(_02412_),
    .C(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__and2_1 _13334_ (.A(_06795_),
    .B(\fifo0.fifo_store[35][7] ),
    .X(_02416_));
 sky130_fd_sc_hd__a211o_1 _13335_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[34][7] ),
    .B1(_02416_),
    .C1(_06728_),
    .X(_02417_));
 sky130_fd_sc_hd__a21o_1 _13336_ (.A1(_07227_),
    .A2(\fifo0.fifo_store[33][7] ),
    .B1(_06528_),
    .X(_02418_));
 sky130_fd_sc_hd__a21o_1 _13337_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[32][7] ),
    .B1(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__a31o_1 _13338_ (.A1(_06681_),
    .A2(_02417_),
    .A3(_02419_),
    .B1(_06630_),
    .X(_02420_));
 sky130_fd_sc_hd__o221a_1 _13339_ (.A1(_02404_),
    .A2(_02410_),
    .B1(_02415_),
    .B2(_02420_),
    .C1(_06679_),
    .X(_02421_));
 sky130_fd_sc_hd__and2_1 _13340_ (.A(_06697_),
    .B(\fifo0.fifo_store[51][7] ),
    .X(_02422_));
 sky130_fd_sc_hd__a211o_1 _13341_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[50][7] ),
    .B1(_02422_),
    .C1(_06650_),
    .X(_02423_));
 sky130_fd_sc_hd__a21o_1 _13342_ (.A1(_06848_),
    .A2(\fifo0.fifo_store[49][7] ),
    .B1(_06725_),
    .X(_02424_));
 sky130_fd_sc_hd__a21o_1 _13343_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[48][7] ),
    .B1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__and2b_1 _13344_ (.A_N(_06586_),
    .B(\fifo0.fifo_store[52][7] ),
    .X(_02426_));
 sky130_fd_sc_hd__a21o_1 _13345_ (.A1(_06536_),
    .A2(\fifo0.fifo_store[53][7] ),
    .B1(_06647_),
    .X(_02427_));
 sky130_fd_sc_hd__and2b_1 _13346_ (.A_N(_06977_),
    .B(\fifo0.fifo_store[54][7] ),
    .X(_02428_));
 sky130_fd_sc_hd__a21bo_1 _13347_ (.A1(_06600_),
    .A2(\fifo0.fifo_store[55][7] ),
    .B1_N(_06420_),
    .X(_02429_));
 sky130_fd_sc_hd__o221a_1 _13348_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_02428_),
    .B2(_02429_),
    .C1(_06655_),
    .X(_02430_));
 sky130_fd_sc_hd__a311o_1 _13349_ (.A1(_06814_),
    .A2(_02423_),
    .A3(_02425_),
    .B1(_06491_),
    .C1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__and2_1 _13350_ (.A(_06697_),
    .B(\fifo0.fifo_store[59][7] ),
    .X(_02432_));
 sky130_fd_sc_hd__a211o_1 _13351_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[58][7] ),
    .B1(_02432_),
    .C1(_06650_),
    .X(_02433_));
 sky130_fd_sc_hd__a21o_1 _13352_ (.A1(_06848_),
    .A2(\fifo0.fifo_store[57][7] ),
    .B1(_06711_),
    .X(_02434_));
 sky130_fd_sc_hd__a21o_1 _13353_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[56][7] ),
    .B1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__and2b_1 _13354_ (.A_N(_06586_),
    .B(\fifo0.fifo_store[62][7] ),
    .X(_02436_));
 sky130_fd_sc_hd__a21bo_1 _13355_ (.A1(_06795_),
    .A2(\fifo0.fifo_store[63][7] ),
    .B1_N(_06578_),
    .X(_02437_));
 sky130_fd_sc_hd__and2b_1 _13356_ (.A_N(_06499_),
    .B(\fifo0.fifo_store[60][7] ),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _13357_ (.A1(_06810_),
    .A2(\fifo0.fifo_store[61][7] ),
    .B1(_06690_),
    .X(_02439_));
 sky130_fd_sc_hd__o221a_1 _13358_ (.A1(_02436_),
    .A2(_02437_),
    .B1(_02438_),
    .B2(_02439_),
    .C1(_06655_),
    .X(_02440_));
 sky130_fd_sc_hd__a311o_1 _13359_ (.A1(_06814_),
    .A2(_02433_),
    .A3(_02435_),
    .B1(_06467_),
    .C1(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__a31o_2 _13360_ (.A1(_06804_),
    .A2(_02431_),
    .A3(_02441_),
    .B1(_06677_),
    .X(_02442_));
 sky130_fd_sc_hd__and2_1 _13361_ (.A(_06499_),
    .B(\fifo0.fifo_store[19][7] ),
    .X(_02443_));
 sky130_fd_sc_hd__a211o_1 _13362_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[18][7] ),
    .B1(_02443_),
    .C1(_06829_),
    .X(_02444_));
 sky130_fd_sc_hd__a21o_1 _13363_ (.A1(_06973_),
    .A2(\fifo0.fifo_store[17][7] ),
    .B1(_07072_),
    .X(_02445_));
 sky130_fd_sc_hd__a21o_1 _13364_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[16][7] ),
    .B1(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__and3_1 _13365_ (.A(_06814_),
    .B(_02444_),
    .C(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__and2_1 _13366_ (.A(_06451_),
    .B(\fifo0.fifo_store[23][7] ),
    .X(_02448_));
 sky130_fd_sc_hd__a211o_1 _13367_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[22][7] ),
    .B1(_02448_),
    .C1(_06728_),
    .X(_02449_));
 sky130_fd_sc_hd__a21o_1 _13368_ (.A1(_06427_),
    .A2(\fifo0.fifo_store[21][7] ),
    .B1(_06975_),
    .X(_02450_));
 sky130_fd_sc_hd__a21o_1 _13369_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[20][7] ),
    .B1(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__a31o_1 _13370_ (.A1(_06824_),
    .A2(_02449_),
    .A3(_02451_),
    .B1(_06630_),
    .X(_02452_));
 sky130_fd_sc_hd__and2_1 _13371_ (.A(_06457_),
    .B(\fifo0.fifo_store[27][7] ),
    .X(_02453_));
 sky130_fd_sc_hd__a211o_1 _13372_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[26][7] ),
    .B1(_02453_),
    .C1(_06728_),
    .X(_02454_));
 sky130_fd_sc_hd__a21o_1 _13373_ (.A1(_06427_),
    .A2(\fifo0.fifo_store[25][7] ),
    .B1(_06975_),
    .X(_02455_));
 sky130_fd_sc_hd__a21o_1 _13374_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[24][7] ),
    .B1(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__and3_1 _13375_ (.A(_06681_),
    .B(_02454_),
    .C(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__a21o_1 _13376_ (.A1(_06959_),
    .A2(\fifo0.fifo_store[29][7] ),
    .B1(_06561_),
    .X(_02458_));
 sky130_fd_sc_hd__a21o_1 _13377_ (.A1(_02205_),
    .A2(\fifo0.fifo_store[28][7] ),
    .B1(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__and2_1 _13378_ (.A(_06521_),
    .B(\fifo0.fifo_store[31][7] ),
    .X(_02460_));
 sky130_fd_sc_hd__a211o_1 _13379_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[30][7] ),
    .B1(_02460_),
    .C1(_06728_),
    .X(_02461_));
 sky130_fd_sc_hd__a31o_1 _13380_ (.A1(_06824_),
    .A2(_02459_),
    .A3(_02461_),
    .B1(_06868_),
    .X(_02462_));
 sky130_fd_sc_hd__o221a_1 _13381_ (.A1(_02447_),
    .A2(_02452_),
    .B1(_02457_),
    .B2(_02462_),
    .C1(_06966_),
    .X(_02463_));
 sky130_fd_sc_hd__and2_1 _13382_ (.A(_02265_),
    .B(\fifo0.fifo_store[11][7] ),
    .X(_02464_));
 sky130_fd_sc_hd__a211o_1 _13383_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[10][7] ),
    .B1(_02464_),
    .C1(_06829_),
    .X(_02465_));
 sky130_fd_sc_hd__a21o_1 _13384_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[9][7] ),
    .B1(_07072_),
    .X(_02466_));
 sky130_fd_sc_hd__a21o_1 _13385_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[8][7] ),
    .B1(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__and2b_1 _13386_ (.A_N(_06591_),
    .B(\fifo0.fifo_store[14][7] ),
    .X(_02468_));
 sky130_fd_sc_hd__a21bo_1 _13387_ (.A1(_06600_),
    .A2(\fifo0.fifo_store[15][7] ),
    .B1_N(_06420_),
    .X(_02469_));
 sky130_fd_sc_hd__and2b_1 _13388_ (.A_N(_06795_),
    .B(\fifo0.fifo_store[12][7] ),
    .X(_02470_));
 sky130_fd_sc_hd__a21o_1 _13389_ (.A1(_07017_),
    .A2(\fifo0.fifo_store[13][7] ),
    .B1(_06984_),
    .X(_02471_));
 sky130_fd_sc_hd__o221a_1 _13390_ (.A1(_02468_),
    .A2(_02469_),
    .B1(_02470_),
    .B2(_02471_),
    .C1(_06683_),
    .X(_02472_));
 sky130_fd_sc_hd__a311o_1 _13391_ (.A1(_06681_),
    .A2(_02465_),
    .A3(_02467_),
    .B1(_06621_),
    .C1(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__and2_1 _13392_ (.A(_02265_),
    .B(\fifo0.fifo_store[3][7] ),
    .X(_02474_));
 sky130_fd_sc_hd__a211o_1 _13393_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[2][7] ),
    .B1(_02474_),
    .C1(_06829_),
    .X(_02475_));
 sky130_fd_sc_hd__a21o_1 _13394_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[1][7] ),
    .B1(_07072_),
    .X(_02476_));
 sky130_fd_sc_hd__a21o_1 _13395_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[0][7] ),
    .B1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__and2b_1 _13396_ (.A_N(_06591_),
    .B(\fifo0.fifo_store[4][7] ),
    .X(_02478_));
 sky130_fd_sc_hd__a21o_1 _13397_ (.A1(_06810_),
    .A2(\fifo0.fifo_store[5][7] ),
    .B1(_06731_),
    .X(_02479_));
 sky130_fd_sc_hd__and2b_1 _13398_ (.A_N(_06795_),
    .B(\fifo0.fifo_store[6][7] ),
    .X(_02480_));
 sky130_fd_sc_hd__a21bo_1 _13399_ (.A1(_07263_),
    .A2(\fifo0.fifo_store[7][7] ),
    .B1_N(_06703_),
    .X(_02481_));
 sky130_fd_sc_hd__o221a_1 _13400_ (.A1(_02478_),
    .A2(_02479_),
    .B1(_02480_),
    .B2(_02481_),
    .C1(_06683_),
    .X(_02482_));
 sky130_fd_sc_hd__a311o_1 _13401_ (.A1(_06681_),
    .A2(_02475_),
    .A3(_02477_),
    .B1(_06491_),
    .C1(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__a31o_1 _13402_ (.A1(_06679_),
    .A2(_02473_),
    .A3(_02483_),
    .B1(_06643_),
    .X(_02484_));
 sky130_fd_sc_hd__o221a_4 _13403_ (.A1(_02421_),
    .A2(_02442_),
    .B1(_02463_),
    .B2(_02484_),
    .C1(_06965_),
    .X(_02485_));
 sky130_fd_sc_hd__a21o_1 _13404_ (.A1(_06956_),
    .A2(\fifo0.fifo_store[109][7] ),
    .B1(_06695_),
    .X(_02486_));
 sky130_fd_sc_hd__a21o_1 _13405_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[108][7] ),
    .B1(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__and2_1 _13406_ (.A(_06586_),
    .B(\fifo0.fifo_store[111][7] ),
    .X(_02488_));
 sky130_fd_sc_hd__a211o_1 _13407_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[110][7] ),
    .B1(_02488_),
    .C1(_06650_),
    .X(_02489_));
 sky130_fd_sc_hd__and2b_1 _13408_ (.A_N(_02265_),
    .B(\fifo0.fifo_store[104][7] ),
    .X(_02490_));
 sky130_fd_sc_hd__a21o_1 _13409_ (.A1(_06521_),
    .A2(\fifo0.fifo_store[105][7] ),
    .B1(_06731_),
    .X(_02491_));
 sky130_fd_sc_hd__and2b_1 _13410_ (.A_N(_06533_),
    .B(\fifo0.fifo_store[106][7] ),
    .X(_02492_));
 sky130_fd_sc_hd__a21bo_1 _13411_ (.A1(_06479_),
    .A2(\fifo0.fifo_store[107][7] ),
    .B1_N(_06614_),
    .X(_02493_));
 sky130_fd_sc_hd__o221a_1 _13412_ (.A1(_02490_),
    .A2(_02491_),
    .B1(_02492_),
    .B2(_02493_),
    .C1(_06668_),
    .X(_02494_));
 sky130_fd_sc_hd__a311o_1 _13413_ (.A1(_06656_),
    .A2(_02487_),
    .A3(_02489_),
    .B1(_06621_),
    .C1(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__and2b_1 _13414_ (.A_N(_06527_),
    .B(\fifo0.fifo_store[100][7] ),
    .X(_02496_));
 sky130_fd_sc_hd__a21o_1 _13415_ (.A1(_02265_),
    .A2(\fifo0.fifo_store[101][7] ),
    .B1(_06614_),
    .X(_02497_));
 sky130_fd_sc_hd__and2b_1 _13416_ (.A_N(_06563_),
    .B(\fifo0.fifo_store[102][7] ),
    .X(_02498_));
 sky130_fd_sc_hd__a21bo_1 _13417_ (.A1(_06533_),
    .A2(\fifo0.fifo_store[103][7] ),
    .B1_N(_06488_),
    .X(_02499_));
 sky130_fd_sc_hd__o221a_1 _13418_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02498_),
    .B2(_02499_),
    .C1(_06623_),
    .X(_02500_));
 sky130_fd_sc_hd__and2b_1 _13419_ (.A_N(_06697_),
    .B(\fifo0.fifo_store[98][7] ),
    .X(_02501_));
 sky130_fd_sc_hd__a21bo_1 _13420_ (.A1(_06533_),
    .A2(\fifo0.fifo_store[99][7] ),
    .B1_N(_06488_),
    .X(_02502_));
 sky130_fd_sc_hd__and2b_1 _13421_ (.A_N(_06469_),
    .B(\fifo0.fifo_store[96][7] ),
    .X(_02503_));
 sky130_fd_sc_hd__a21o_1 _13422_ (.A1(_06521_),
    .A2(\fifo0.fifo_store[97][7] ),
    .B1(_06731_),
    .X(_02504_));
 sky130_fd_sc_hd__o221a_1 _13423_ (.A1(_02501_),
    .A2(_02502_),
    .B1(_02503_),
    .B2(_02504_),
    .C1(_06634_),
    .X(_02505_));
 sky130_fd_sc_hd__o31a_1 _13424_ (.A1(_06571_),
    .A2(_02500_),
    .A3(_02505_),
    .B1(_06493_),
    .X(_02506_));
 sky130_fd_sc_hd__and2_1 _13425_ (.A(_02265_),
    .B(\fifo0.fifo_store[115][7] ),
    .X(_02507_));
 sky130_fd_sc_hd__a211o_1 _13426_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[114][7] ),
    .B1(_02507_),
    .C1(_06829_),
    .X(_02508_));
 sky130_fd_sc_hd__a21o_1 _13427_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[113][7] ),
    .B1(_06695_),
    .X(_02509_));
 sky130_fd_sc_hd__a21o_1 _13428_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[112][7] ),
    .B1(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__and2b_1 _13429_ (.A_N(_06591_),
    .B(\fifo0.fifo_store[116][7] ),
    .X(_02511_));
 sky130_fd_sc_hd__a21o_1 _13430_ (.A1(_06810_),
    .A2(\fifo0.fifo_store[117][7] ),
    .B1(_06731_),
    .X(_02512_));
 sky130_fd_sc_hd__and2b_1 _13431_ (.A_N(_06795_),
    .B(\fifo0.fifo_store[118][7] ),
    .X(_02513_));
 sky130_fd_sc_hd__a21bo_1 _13432_ (.A1(_07263_),
    .A2(\fifo0.fifo_store[119][7] ),
    .B1_N(_06703_),
    .X(_02514_));
 sky130_fd_sc_hd__o221a_1 _13433_ (.A1(_02511_),
    .A2(_02512_),
    .B1(_02513_),
    .B2(_02514_),
    .C1(_06683_),
    .X(_02515_));
 sky130_fd_sc_hd__a311o_1 _13434_ (.A1(_06681_),
    .A2(_02508_),
    .A3(_02510_),
    .B1(_06491_),
    .C1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__and2b_1 _13435_ (.A_N(_06563_),
    .B(\fifo0.fifo_store[122][7] ),
    .X(_02517_));
 sky130_fd_sc_hd__a21bo_1 _13436_ (.A1(_06499_),
    .A2(\fifo0.fifo_store[123][7] ),
    .B1_N(_06480_),
    .X(_02518_));
 sky130_fd_sc_hd__and2b_1 _13437_ (.A_N(_06697_),
    .B(\fifo0.fifo_store[120][7] ),
    .X(_02519_));
 sky130_fd_sc_hd__a21o_1 _13438_ (.A1(_06503_),
    .A2(\fifo0.fifo_store[121][7] ),
    .B1(_06647_),
    .X(_02520_));
 sky130_fd_sc_hd__o221a_1 _13439_ (.A1(_02517_),
    .A2(_02518_),
    .B1(_02519_),
    .B2(_02520_),
    .C1(_06660_),
    .X(_02521_));
 sky130_fd_sc_hd__and2b_1 _13440_ (.A_N(_06586_),
    .B(\fifo0.fifo_store[124][7] ),
    .X(_02522_));
 sky130_fd_sc_hd__a21o_1 _13441_ (.A1(_06536_),
    .A2(\fifo0.fifo_store[125][7] ),
    .B1(_06647_),
    .X(_02523_));
 sky130_fd_sc_hd__and2b_1 _13442_ (.A_N(_06977_),
    .B(\fifo0.fifo_store[126][7] ),
    .X(_02524_));
 sky130_fd_sc_hd__a21bo_1 _13443_ (.A1(_06600_),
    .A2(\fifo0.fifo_store[127][7] ),
    .B1_N(_06420_),
    .X(_02525_));
 sky130_fd_sc_hd__o221a_1 _13444_ (.A1(_02522_),
    .A2(_02523_),
    .B1(_02524_),
    .B2(_02525_),
    .C1(_06655_),
    .X(_02526_));
 sky130_fd_sc_hd__o31a_1 _13445_ (.A1(_06467_),
    .A2(_02521_),
    .A3(_02526_),
    .B1(_06641_),
    .X(_02527_));
 sky130_fd_sc_hd__a221o_4 _13446_ (.A1(_02495_),
    .A2(_02506_),
    .B1(_02516_),
    .B2(_02527_),
    .C1(_06677_),
    .X(_02528_));
 sky130_fd_sc_hd__and2_1 _13447_ (.A(_06586_),
    .B(\fifo0.fifo_store[83][7] ),
    .X(_02529_));
 sky130_fd_sc_hd__a211o_1 _13448_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[82][7] ),
    .B1(_02529_),
    .C1(_06650_),
    .X(_02530_));
 sky130_fd_sc_hd__a21o_1 _13449_ (.A1(_06658_),
    .A2(\fifo0.fifo_store[81][7] ),
    .B1(_06725_),
    .X(_02531_));
 sky130_fd_sc_hd__a21o_1 _13450_ (.A1(_06993_),
    .A2(\fifo0.fifo_store[80][7] ),
    .B1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__and2b_1 _13451_ (.A_N(_06469_),
    .B(\fifo0.fifo_store[84][7] ),
    .X(_02533_));
 sky130_fd_sc_hd__a21o_1 _13452_ (.A1(_06521_),
    .A2(\fifo0.fifo_store[85][7] ),
    .B1(_06647_),
    .X(_02534_));
 sky130_fd_sc_hd__and2b_1 _13453_ (.A_N(_06591_),
    .B(\fifo0.fifo_store[86][7] ),
    .X(_02535_));
 sky130_fd_sc_hd__a21bo_1 _13454_ (.A1(_06810_),
    .A2(\fifo0.fifo_store[87][7] ),
    .B1_N(_06420_),
    .X(_02536_));
 sky130_fd_sc_hd__o221a_2 _13455_ (.A1(_02533_),
    .A2(_02534_),
    .B1(_02535_),
    .B2(_02536_),
    .C1(_06655_),
    .X(_02537_));
 sky130_fd_sc_hd__a311o_1 _13456_ (.A1(_06814_),
    .A2(_02530_),
    .A3(_02532_),
    .B1(_06491_),
    .C1(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__and2b_1 _13457_ (.A_N(_06527_),
    .B(\fifo0.fifo_store[90][7] ),
    .X(_02539_));
 sky130_fd_sc_hd__a21bo_1 _13458_ (.A1(_06469_),
    .A2(\fifo0.fifo_store[91][7] ),
    .B1_N(_06627_),
    .X(_02540_));
 sky130_fd_sc_hd__and2b_1 _13459_ (.A_N(_06563_),
    .B(\fifo0.fifo_store[88][7] ),
    .X(_02541_));
 sky130_fd_sc_hd__a21o_1 _13460_ (.A1(_06457_),
    .A2(\fifo0.fifo_store[89][7] ),
    .B1(_06718_),
    .X(_02542_));
 sky130_fd_sc_hd__o221a_1 _13461_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02541_),
    .B2(_02542_),
    .C1(_06660_),
    .X(_02543_));
 sky130_fd_sc_hd__and2b_1 _13462_ (.A_N(_06434_),
    .B(\fifo0.fifo_store[92][7] ),
    .X(_02544_));
 sky130_fd_sc_hd__a21o_1 _13463_ (.A1(_06451_),
    .A2(\fifo0.fifo_store[93][7] ),
    .B1(_06718_),
    .X(_02545_));
 sky130_fd_sc_hd__and2b_1 _13464_ (.A_N(_06469_),
    .B(\fifo0.fifo_store[94][7] ),
    .X(_02546_));
 sky130_fd_sc_hd__a21bo_1 _13465_ (.A1(_06536_),
    .A2(\fifo0.fifo_store[95][7] ),
    .B1_N(_06510_),
    .X(_02547_));
 sky130_fd_sc_hd__o221a_1 _13466_ (.A1(_02544_),
    .A2(_02545_),
    .B1(_02546_),
    .B2(_02547_),
    .C1(_06655_),
    .X(_02548_));
 sky130_fd_sc_hd__o31a_1 _13467_ (.A1(_06467_),
    .A2(_02543_),
    .A3(_02548_),
    .B1(_06641_),
    .X(_02549_));
 sky130_fd_sc_hd__a21o_1 _13468_ (.A1(_06801_),
    .A2(\fifo0.fifo_store[77][7] ),
    .B1(_07072_),
    .X(_02550_));
 sky130_fd_sc_hd__a21o_1 _13469_ (.A1(_07077_),
    .A2(\fifo0.fifo_store[76][7] ),
    .B1(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__and2_1 _13470_ (.A(_02265_),
    .B(\fifo0.fifo_store[79][7] ),
    .X(_02552_));
 sky130_fd_sc_hd__a211o_1 _13471_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[78][7] ),
    .B1(_02552_),
    .C1(_06829_),
    .X(_02553_));
 sky130_fd_sc_hd__and2b_1 _13472_ (.A_N(_06977_),
    .B(\fifo0.fifo_store[72][7] ),
    .X(_02554_));
 sky130_fd_sc_hd__a21o_1 _13473_ (.A1(_06810_),
    .A2(\fifo0.fifo_store[73][7] ),
    .B1(_06731_),
    .X(_02555_));
 sky130_fd_sc_hd__and2b_1 _13474_ (.A_N(_06451_),
    .B(\fifo0.fifo_store[74][7] ),
    .X(_02556_));
 sky130_fd_sc_hd__a21bo_1 _13475_ (.A1(_07263_),
    .A2(\fifo0.fifo_store[75][7] ),
    .B1_N(_06703_),
    .X(_02557_));
 sky130_fd_sc_hd__o221a_1 _13476_ (.A1(_02554_),
    .A2(_02555_),
    .B1(_02556_),
    .B2(_02557_),
    .C1(_06668_),
    .X(_02558_));
 sky130_fd_sc_hd__a311o_1 _13477_ (.A1(_06656_),
    .A2(_02551_),
    .A3(_02553_),
    .B1(_06621_),
    .C1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__and2b_1 _13478_ (.A_N(_06563_),
    .B(\fifo0.fifo_store[68][7] ),
    .X(_02560_));
 sky130_fd_sc_hd__a21o_1 _13479_ (.A1(_06591_),
    .A2(\fifo0.fifo_store[69][7] ),
    .B1(_06718_),
    .X(_02561_));
 sky130_fd_sc_hd__and2b_1 _13480_ (.A_N(_06697_),
    .B(\fifo0.fifo_store[70][7] ),
    .X(_02562_));
 sky130_fd_sc_hd__a21bo_1 _13481_ (.A1(_06451_),
    .A2(\fifo0.fifo_store[71][7] ),
    .B1_N(_06578_),
    .X(_02563_));
 sky130_fd_sc_hd__o221a_1 _13482_ (.A1(_02560_),
    .A2(_02561_),
    .B1(_02562_),
    .B2(_02563_),
    .C1(_06623_),
    .X(_02564_));
 sky130_fd_sc_hd__and2b_1 _13483_ (.A_N(_06586_),
    .B(\fifo0.fifo_store[66][7] ),
    .X(_02565_));
 sky130_fd_sc_hd__a21bo_1 _13484_ (.A1(_06795_),
    .A2(\fifo0.fifo_store[67][7] ),
    .B1_N(_06578_),
    .X(_02566_));
 sky130_fd_sc_hd__and2b_1 _13485_ (.A_N(_06499_),
    .B(\fifo0.fifo_store[64][7] ),
    .X(_02567_));
 sky130_fd_sc_hd__a21o_1 _13486_ (.A1(_06479_),
    .A2(\fifo0.fifo_store[65][7] ),
    .B1(_06690_),
    .X(_02568_));
 sky130_fd_sc_hd__o221a_1 _13487_ (.A1(_02565_),
    .A2(_02566_),
    .B1(_02567_),
    .B2(_02568_),
    .C1(_06668_),
    .X(_02569_));
 sky130_fd_sc_hd__o31a_1 _13488_ (.A1(_06491_),
    .A2(_02564_),
    .A3(_02569_),
    .B1(_06743_),
    .X(_02570_));
 sky130_fd_sc_hd__a221o_2 _13489_ (.A1(_02538_),
    .A2(_02549_),
    .B1(_02559_),
    .B2(_02570_),
    .C1(_00005_),
    .X(_02571_));
 sky130_fd_sc_hd__a31o_2 _13490_ (.A1(_06992_),
    .A2(_02528_),
    .A3(_02571_),
    .B1(net23),
    .X(_02572_));
 sky130_fd_sc_hd__o32a_2 _13491_ (.A1(_06357_),
    .A2(_02393_),
    .A3(_02398_),
    .B1(_02485_),
    .B2(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(_02370_),
    .A1(_02573_),
    .S(_07164_),
    .X(_02574_));
 sky130_fd_sc_hd__mux4_1 _13493_ (.A0(\fifo0.fifo_store[36][5] ),
    .A1(\fifo0.fifo_store[37][5] ),
    .A2(\fifo0.fifo_store[38][5] ),
    .A3(\fifo0.fifo_store[39][5] ),
    .S0(_06625_),
    .S1(_06489_),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_1 _13494_ (.A0(\fifo0.fifo_store[32][5] ),
    .A1(\fifo0.fifo_store[33][5] ),
    .A2(\fifo0.fifo_store[34][5] ),
    .A3(\fifo0.fifo_store[35][5] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_02576_));
 sky130_fd_sc_hd__or2_1 _13495_ (.A(_06484_),
    .B(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__o211a_1 _13496_ (.A1(_07371_),
    .A2(_02575_),
    .B1(_02577_),
    .C1(_06868_),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_1 _13497_ (.A0(\fifo0.fifo_store[40][5] ),
    .A1(\fifo0.fifo_store[41][5] ),
    .A2(\fifo0.fifo_store[42][5] ),
    .A3(\fifo0.fifo_store[43][5] ),
    .S0(_06956_),
    .S1(_06421_),
    .X(_02579_));
 sky130_fd_sc_hd__or2b_1 _13498_ (.A(\fifo0.fifo_store[47][5] ),
    .B_N(_06533_),
    .X(_02580_));
 sky130_fd_sc_hd__o21a_1 _13499_ (.A1(_06533_),
    .A2(\fifo0.fifo_store[46][5] ),
    .B1(_06647_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(\fifo0.fifo_store[44][5] ),
    .A1(\fifo0.fifo_store[45][5] ),
    .S(_06710_),
    .X(_02582_));
 sky130_fd_sc_hd__a221o_1 _13501_ (.A1(_02580_),
    .A2(_02581_),
    .B1(_02582_),
    .B2(_06650_),
    .C1(_06660_),
    .X(_02583_));
 sky130_fd_sc_hd__o211a_1 _13502_ (.A1(_06656_),
    .A2(_02579_),
    .B1(_02583_),
    .C1(_06664_),
    .X(_02584_));
 sky130_fd_sc_hd__mux4_1 _13503_ (.A0(\fifo0.fifo_store[48][5] ),
    .A1(\fifo0.fifo_store[49][5] ),
    .A2(\fifo0.fifo_store[50][5] ),
    .A3(\fifo0.fifo_store[51][5] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_02585_));
 sky130_fd_sc_hd__mux4_1 _13504_ (.A0(\fifo0.fifo_store[52][5] ),
    .A1(\fifo0.fifo_store[53][5] ),
    .A2(\fifo0.fifo_store[54][5] ),
    .A3(\fifo0.fifo_store[55][5] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(_02585_),
    .A1(_02586_),
    .S(_06440_),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_1 _13506_ (.A0(\fifo0.fifo_store[60][5] ),
    .A1(\fifo0.fifo_store[61][5] ),
    .A2(\fifo0.fifo_store[62][5] ),
    .A3(\fifo0.fifo_store[63][5] ),
    .S0(_06673_),
    .S1(_06420_),
    .X(_02588_));
 sky130_fd_sc_hd__or2_1 _13507_ (.A(_06668_),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__mux4_1 _13508_ (.A0(\fifo0.fifo_store[56][5] ),
    .A1(\fifo0.fifo_store[57][5] ),
    .A2(\fifo0.fifo_store[58][5] ),
    .A3(\fifo0.fifo_store[59][5] ),
    .S0(_06717_),
    .S1(_06718_),
    .X(_02590_));
 sky130_fd_sc_hd__o21a_1 _13509_ (.A1(_06730_),
    .A2(_02590_),
    .B1(_06663_),
    .X(_02591_));
 sky130_fd_sc_hd__a221o_2 _13510_ (.A1(_06735_),
    .A2(_02587_),
    .B1(_02589_),
    .B2(_02591_),
    .C1(_06743_),
    .X(_02592_));
 sky130_fd_sc_hd__o311a_1 _13511_ (.A1(_06589_),
    .A2(_02578_),
    .A3(_02584_),
    .B1(_06643_),
    .C1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__mux4_1 _13512_ (.A0(\fifo0.fifo_store[28][5] ),
    .A1(\fifo0.fifo_store[29][5] ),
    .A2(\fifo0.fifo_store[30][5] ),
    .A3(\fifo0.fifo_store[31][5] ),
    .S0(_06848_),
    .S1(_06579_),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_2 _13513_ (.A0(\fifo0.fifo_store[24][5] ),
    .A1(\fifo0.fifo_store[25][5] ),
    .A2(\fifo0.fifo_store[26][5] ),
    .A3(\fifo0.fifo_store[27][5] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_02595_));
 sky130_fd_sc_hd__or2_1 _13514_ (.A(_06484_),
    .B(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__o211a_1 _13515_ (.A1(_06814_),
    .A2(_02594_),
    .B1(_02596_),
    .C1(_06630_),
    .X(_02597_));
 sky130_fd_sc_hd__or2_1 _13516_ (.A(_06499_),
    .B(\fifo0.fifo_store[20][5] ),
    .X(_02598_));
 sky130_fd_sc_hd__o211a_1 _13517_ (.A1(_02399_),
    .A2(\fifo0.fifo_store[21][5] ),
    .B1(_02598_),
    .C1(_06728_),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(\fifo0.fifo_store[22][5] ),
    .A1(\fifo0.fifo_store[23][5] ),
    .S(_06544_),
    .X(_02600_));
 sky130_fd_sc_hd__a21o_1 _13519_ (.A1(_06971_),
    .A2(_02600_),
    .B1(_06634_),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_2 _13520_ (.A0(\fifo0.fifo_store[16][5] ),
    .A1(\fifo0.fifo_store[17][5] ),
    .A2(\fifo0.fifo_store[18][5] ),
    .A3(\fifo0.fifo_store[19][5] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_02602_));
 sky130_fd_sc_hd__o221a_1 _13521_ (.A1(_02599_),
    .A2(_02601_),
    .B1(_02602_),
    .B2(_06656_),
    .C1(_06735_),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_1 _13522_ (.A0(\fifo0.fifo_store[12][5] ),
    .A1(\fifo0.fifo_store[13][5] ),
    .A2(\fifo0.fifo_store[14][5] ),
    .A3(\fifo0.fifo_store[15][5] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_02604_));
 sky130_fd_sc_hd__or2_1 _13523_ (.A(_06634_),
    .B(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__mux4_2 _13524_ (.A0(\fifo0.fifo_store[8][5] ),
    .A1(\fifo0.fifo_store[9][5] ),
    .A2(\fifo0.fifo_store[10][5] ),
    .A3(\fifo0.fifo_store[11][5] ),
    .S0(_06548_),
    .S1(_06614_),
    .X(_02606_));
 sky130_fd_sc_hd__o21a_1 _13525_ (.A1(_06683_),
    .A2(_02606_),
    .B1(_06663_),
    .X(_02607_));
 sky130_fd_sc_hd__mux4_1 _13526_ (.A0(\fifo0.fifo_store[4][5] ),
    .A1(\fifo0.fifo_store[5][5] ),
    .A2(\fifo0.fifo_store[6][5] ),
    .A3(\fifo0.fifo_store[7][5] ),
    .S0(_06673_),
    .S1(_06510_),
    .X(_02608_));
 sky130_fd_sc_hd__or2_1 _13527_ (.A(_06668_),
    .B(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__mux4_1 _13528_ (.A0(\fifo0.fifo_store[0][5] ),
    .A1(\fifo0.fifo_store[1][5] ),
    .A2(\fifo0.fifo_store[2][5] ),
    .A3(\fifo0.fifo_store[3][5] ),
    .S0(_06717_),
    .S1(_06703_),
    .X(_02610_));
 sky130_fd_sc_hd__o21a_1 _13529_ (.A1(_06730_),
    .A2(_02610_),
    .B1(_06466_),
    .X(_02611_));
 sky130_fd_sc_hd__a221o_1 _13530_ (.A1(_02605_),
    .A2(_02607_),
    .B1(_02609_),
    .B2(_02611_),
    .C1(_06641_),
    .X(_02612_));
 sky130_fd_sc_hd__o311a_1 _13531_ (.A1(_06679_),
    .A2(_02597_),
    .A3(_02603_),
    .B1(_02612_),
    .C1(_06677_),
    .X(_02613_));
 sky130_fd_sc_hd__or3_4 _13532_ (.A(_00006_),
    .B(_02593_),
    .C(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_1 _13533_ (.A0(\fifo0.fifo_store[100][5] ),
    .A1(\fifo0.fifo_store[101][5] ),
    .A2(\fifo0.fifo_store[102][5] ),
    .A3(\fifo0.fifo_store[103][5] ),
    .S0(_06693_),
    .S1(_06579_),
    .X(_02615_));
 sky130_fd_sc_hd__mux4_1 _13534_ (.A0(\fifo0.fifo_store[96][5] ),
    .A1(\fifo0.fifo_store[97][5] ),
    .A2(\fifo0.fifo_store[98][5] ),
    .A3(\fifo0.fifo_store[99][5] ),
    .S0(_06486_),
    .S1(_06480_),
    .X(_02616_));
 sky130_fd_sc_hd__or2_1 _13535_ (.A(_06484_),
    .B(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__o211a_1 _13536_ (.A1(_06814_),
    .A2(_02615_),
    .B1(_02617_),
    .C1(_06868_),
    .X(_02618_));
 sky130_fd_sc_hd__mux4_2 _13537_ (.A0(\fifo0.fifo_store[104][5] ),
    .A1(\fifo0.fifo_store[105][5] ),
    .A2(\fifo0.fifo_store[106][5] ),
    .A3(\fifo0.fifo_store[107][5] ),
    .S0(_06973_),
    .S1(_06421_),
    .X(_02619_));
 sky130_fd_sc_hd__or2b_1 _13538_ (.A(\fifo0.fifo_store[111][5] ),
    .B_N(_06503_),
    .X(_02620_));
 sky130_fd_sc_hd__o21a_1 _13539_ (.A1(_06503_),
    .A2(\fifo0.fifo_store[110][5] ),
    .B1(_06731_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(\fifo0.fifo_store[108][5] ),
    .A1(\fifo0.fifo_store[109][5] ),
    .S(_07008_),
    .X(_02622_));
 sky130_fd_sc_hd__a221o_1 _13541_ (.A1(_02620_),
    .A2(_02621_),
    .B1(_02622_),
    .B2(_06829_),
    .C1(_06634_),
    .X(_02623_));
 sky130_fd_sc_hd__o211a_1 _13542_ (.A1(_06656_),
    .A2(_02619_),
    .B1(_02623_),
    .C1(_06664_),
    .X(_02624_));
 sky130_fd_sc_hd__mux4_1 _13543_ (.A0(\fifo0.fifo_store[112][5] ),
    .A1(\fifo0.fifo_store[113][5] ),
    .A2(\fifo0.fifo_store[114][5] ),
    .A3(\fifo0.fifo_store[115][5] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_1 _13544_ (.A0(\fifo0.fifo_store[116][5] ),
    .A1(\fifo0.fifo_store[117][5] ),
    .A2(\fifo0.fifo_store[118][5] ),
    .A3(\fifo0.fifo_store[119][5] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(_02625_),
    .A1(_02626_),
    .S(_06440_),
    .X(_02627_));
 sky130_fd_sc_hd__mux4_1 _13546_ (.A0(\fifo0.fifo_store[124][5] ),
    .A1(\fifo0.fifo_store[125][5] ),
    .A2(\fifo0.fifo_store[126][5] ),
    .A3(\fifo0.fifo_store[127][5] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_02628_));
 sky130_fd_sc_hd__or2_1 _13547_ (.A(_06634_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__mux4_2 _13548_ (.A0(\fifo0.fifo_store[120][5] ),
    .A1(\fifo0.fifo_store[121][5] ),
    .A2(\fifo0.fifo_store[122][5] ),
    .A3(\fifo0.fifo_store[123][5] ),
    .S0(_06548_),
    .S1(_06703_),
    .X(_02630_));
 sky130_fd_sc_hd__o21a_1 _13549_ (.A1(_06683_),
    .A2(_02630_),
    .B1(_06663_),
    .X(_02631_));
 sky130_fd_sc_hd__a221o_1 _13550_ (.A1(_06868_),
    .A2(_02627_),
    .B1(_02629_),
    .B2(_02631_),
    .C1(_06743_),
    .X(_02632_));
 sky130_fd_sc_hd__o311a_1 _13551_ (.A1(_06804_),
    .A2(_02618_),
    .A3(_02624_),
    .B1(_02632_),
    .C1(_06643_),
    .X(_02633_));
 sky130_fd_sc_hd__mux4_1 _13552_ (.A0(\fifo0.fifo_store[76][5] ),
    .A1(\fifo0.fifo_store[77][5] ),
    .A2(\fifo0.fifo_store[78][5] ),
    .A3(\fifo0.fifo_store[79][5] ),
    .S0(_06956_),
    .S1(_06421_),
    .X(_02634_));
 sky130_fd_sc_hd__mux4_1 _13553_ (.A0(\fifo0.fifo_store[72][5] ),
    .A1(\fifo0.fifo_store[73][5] ),
    .A2(\fifo0.fifo_store[74][5] ),
    .A3(\fifo0.fifo_store[75][5] ),
    .S0(_06426_),
    .S1(_06488_),
    .X(_02635_));
 sky130_fd_sc_hd__or2_1 _13554_ (.A(_06623_),
    .B(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__o211a_1 _13555_ (.A1(_06814_),
    .A2(_02634_),
    .B1(_02636_),
    .C1(_06664_),
    .X(_02637_));
 sky130_fd_sc_hd__or2_1 _13556_ (.A(_06533_),
    .B(\fifo0.fifo_store[68][5] ),
    .X(_02638_));
 sky130_fd_sc_hd__o211a_1 _13557_ (.A1(_02407_),
    .A2(\fifo0.fifo_store[69][5] ),
    .B1(_02638_),
    .C1(_06728_),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(\fifo0.fifo_store[70][5] ),
    .A1(\fifo0.fifo_store[71][5] ),
    .S(_06507_),
    .X(_02640_));
 sky130_fd_sc_hd__a21o_1 _13559_ (.A1(_06971_),
    .A2(_02640_),
    .B1(_06668_),
    .X(_02641_));
 sky130_fd_sc_hd__mux4_1 _13560_ (.A0(\fifo0.fifo_store[64][5] ),
    .A1(\fifo0.fifo_store[65][5] ),
    .A2(\fifo0.fifo_store[66][5] ),
    .A3(\fifo0.fifo_store[67][5] ),
    .S0(_06973_),
    .S1(_06421_),
    .X(_02642_));
 sky130_fd_sc_hd__o221a_1 _13561_ (.A1(_02639_),
    .A2(_02641_),
    .B1(_02642_),
    .B2(_06824_),
    .C1(_06735_),
    .X(_02643_));
 sky130_fd_sc_hd__mux4_1 _13562_ (.A0(\fifo0.fifo_store[88][5] ),
    .A1(\fifo0.fifo_store[89][5] ),
    .A2(\fifo0.fifo_store[90][5] ),
    .A3(\fifo0.fifo_store[91][5] ),
    .S0(_06673_),
    .S1(_06420_),
    .X(_02644_));
 sky130_fd_sc_hd__or2_1 _13563_ (.A(_06655_),
    .B(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_2 _13564_ (.A0(\fifo0.fifo_store[92][5] ),
    .A1(\fifo0.fifo_store[93][5] ),
    .A2(\fifo0.fifo_store[94][5] ),
    .A3(\fifo0.fifo_store[95][5] ),
    .S0(_06717_),
    .S1(_06718_),
    .X(_02646_));
 sky130_fd_sc_hd__o21a_1 _13565_ (.A1(_06680_),
    .A2(_02646_),
    .B1(_06663_),
    .X(_02647_));
 sky130_fd_sc_hd__mux4_1 _13566_ (.A0(\fifo0.fifo_store[84][5] ),
    .A1(\fifo0.fifo_store[85][5] ),
    .A2(\fifo0.fifo_store[86][5] ),
    .A3(\fifo0.fifo_store[87][5] ),
    .S0(_06548_),
    .S1(_06614_),
    .X(_02648_));
 sky130_fd_sc_hd__or2_1 _13567_ (.A(_06668_),
    .B(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__mux4_1 _13568_ (.A0(\fifo0.fifo_store[80][5] ),
    .A1(\fifo0.fifo_store[81][5] ),
    .A2(\fifo0.fifo_store[82][5] ),
    .A3(\fifo0.fifo_store[83][5] ),
    .S0(_06513_),
    .S1(_06718_),
    .X(_02650_));
 sky130_fd_sc_hd__o21a_1 _13569_ (.A1(_06730_),
    .A2(_02650_),
    .B1(_06466_),
    .X(_02651_));
 sky130_fd_sc_hd__a221o_1 _13570_ (.A1(_02645_),
    .A2(_02647_),
    .B1(_02649_),
    .B2(_02651_),
    .C1(_06743_),
    .X(_02652_));
 sky130_fd_sc_hd__o311a_1 _13571_ (.A1(_06804_),
    .A2(_02637_),
    .A3(_02643_),
    .B1(_02652_),
    .C1(_06677_),
    .X(_02653_));
 sky130_fd_sc_hd__or3_4 _13572_ (.A(_06965_),
    .B(_02633_),
    .C(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__and2_1 _13573_ (.A(_06753_),
    .B(_06778_),
    .X(_02655_));
 sky130_fd_sc_hd__a21oi_1 _13574_ (.A1(_06892_),
    .A2(_07421_),
    .B1(_06396_),
    .Y(_02656_));
 sky130_fd_sc_hd__a31o_1 _13575_ (.A1(_06363_),
    .A2(_06897_),
    .A3(_06905_),
    .B1(_06358_),
    .X(_02657_));
 sky130_fd_sc_hd__o311a_1 _13576_ (.A1(_06402_),
    .A2(_02655_),
    .A3(_02656_),
    .B1(_02657_),
    .C1(_06404_),
    .X(_02658_));
 sky130_fd_sc_hd__nor2_1 _13577_ (.A(_06751_),
    .B(_06775_),
    .Y(_02659_));
 sky130_fd_sc_hd__o21ai_1 _13578_ (.A1(_07042_),
    .A2(_06781_),
    .B1(_06786_),
    .Y(_02660_));
 sky130_fd_sc_hd__o21a_1 _13579_ (.A1(_02659_),
    .A2(_02660_),
    .B1(_07193_),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _13580_ (.A(_06922_),
    .B(_06759_),
    .Y(_02662_));
 sky130_fd_sc_hd__and4_1 _13581_ (.A(_06764_),
    .B(_06766_),
    .C(_06910_),
    .D(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__o31ai_1 _13582_ (.A1(_02658_),
    .A2(_02661_),
    .A3(_02663_),
    .B1(_06769_),
    .Y(_02664_));
 sky130_fd_sc_hd__and2_1 _13583_ (.A(_07193_),
    .B(_06400_),
    .X(_02665_));
 sky130_fd_sc_hd__nor2_1 _13584_ (.A(_06747_),
    .B(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__o41a_1 _13585_ (.A1(_02658_),
    .A2(_02661_),
    .A3(_02663_),
    .A4(_02666_),
    .B1(_06918_),
    .X(_02667_));
 sky130_fd_sc_hd__a32o_1 _13586_ (.A1(_06606_),
    .A2(_02614_),
    .A3(_02654_),
    .B1(_02664_),
    .B2(_02667_),
    .X(_02668_));
 sky130_fd_sc_hd__mux4_1 _13587_ (.A0(\fifo0.fifo_store[96][6] ),
    .A1(\fifo0.fifo_store[97][6] ),
    .A2(\fifo0.fifo_store[98][6] ),
    .A3(\fifo0.fifo_store[99][6] ),
    .S0(_06451_),
    .S1(_06453_),
    .X(_02669_));
 sky130_fd_sc_hd__or2_1 _13588_ (.A(_06448_),
    .B(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__mux4_1 _13589_ (.A0(\fifo0.fifo_store[100][6] ),
    .A1(\fifo0.fifo_store[101][6] ),
    .A2(\fifo0.fifo_store[102][6] ),
    .A3(\fifo0.fifo_store[103][6] ),
    .S0(_06451_),
    .S1(_06453_),
    .X(_02671_));
 sky130_fd_sc_hd__or2_1 _13590_ (.A(_06456_),
    .B(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__mux4_1 _13591_ (.A0(\fifo0.fifo_store[108][6] ),
    .A1(\fifo0.fifo_store[109][6] ),
    .A2(\fifo0.fifo_store[110][6] ),
    .A3(\fifo0.fifo_store[111][6] ),
    .S0(_07017_),
    .S1(_07391_),
    .X(_02673_));
 sky130_fd_sc_hd__mux4_2 _13592_ (.A0(\fifo0.fifo_store[104][6] ),
    .A1(\fifo0.fifo_store[105][6] ),
    .A2(\fifo0.fifo_store[106][6] ),
    .A3(\fifo0.fifo_store[107][6] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02674_));
 sky130_fd_sc_hd__or2_1 _13593_ (.A(_06447_),
    .B(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__o211a_1 _13594_ (.A1(_07371_),
    .A2(_02673_),
    .B1(_02675_),
    .C1(_07219_),
    .X(_02676_));
 sky130_fd_sc_hd__a311o_1 _13595_ (.A1(_06468_),
    .A2(_02670_),
    .A3(_02672_),
    .B1(_06589_),
    .C1(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__or2_1 _13596_ (.A(_06612_),
    .B(\fifo0.fifo_store[127][6] ),
    .X(_02678_));
 sky130_fd_sc_hd__o21a_1 _13597_ (.A1(_07097_),
    .A2(\fifo0.fifo_store[126][6] ),
    .B1(_06615_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(\fifo0.fifo_store[124][6] ),
    .A1(\fifo0.fifo_store[125][6] ),
    .S(_06689_),
    .X(_02680_));
 sky130_fd_sc_hd__a221o_1 _13599_ (.A1(_02678_),
    .A2(_02679_),
    .B1(_02680_),
    .B2(_06425_),
    .C1(_06477_),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_2 _13600_ (.A0(\fifo0.fifo_store[120][6] ),
    .A1(\fifo0.fifo_store[121][6] ),
    .A2(\fifo0.fifo_store[122][6] ),
    .A3(\fifo0.fifo_store[123][6] ),
    .S0(_07263_),
    .S1(_07391_),
    .X(_02682_));
 sky130_fd_sc_hd__o21a_1 _13601_ (.A1(_06485_),
    .A2(_02682_),
    .B1(_06491_),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_1 _13602_ (.A0(\fifo0.fifo_store[112][6] ),
    .A1(\fifo0.fifo_store[113][6] ),
    .A2(\fifo0.fifo_store[114][6] ),
    .A3(\fifo0.fifo_store[115][6] ),
    .S0(_06795_),
    .S1(_06453_),
    .X(_02684_));
 sky130_fd_sc_hd__mux4_1 _13603_ (.A0(\fifo0.fifo_store[116][6] ),
    .A1(\fifo0.fifo_store[117][6] ),
    .A2(\fifo0.fifo_store[118][6] ),
    .A3(\fifo0.fifo_store[119][6] ),
    .S0(_06451_),
    .S1(_06453_),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _13604_ (.A0(_02684_),
    .A1(_02685_),
    .S(_06797_),
    .X(_02686_));
 sky130_fd_sc_hd__a221o_1 _13605_ (.A1(_02681_),
    .A2(_02683_),
    .B1(_02686_),
    .B2(_06468_),
    .C1(_06494_),
    .X(_02687_));
 sky130_fd_sc_hd__or2_1 _13606_ (.A(_06507_),
    .B(\fifo0.fifo_store[94][6] ),
    .X(_02688_));
 sky130_fd_sc_hd__o211a_1 _13607_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[95][6] ),
    .B1(_02688_),
    .C1(_06648_),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_1 _13608_ (.A0(\fifo0.fifo_store[92][6] ),
    .A1(\fifo0.fifo_store[93][6] ),
    .S(_06617_),
    .X(_02690_));
 sky130_fd_sc_hd__a21o_1 _13609_ (.A1(_06650_),
    .A2(_02690_),
    .B1(_06476_),
    .X(_02691_));
 sky130_fd_sc_hd__mux4_2 _13610_ (.A0(\fifo0.fifo_store[88][6] ),
    .A1(\fifo0.fifo_store[89][6] ),
    .A2(\fifo0.fifo_store[90][6] ),
    .A3(\fifo0.fifo_store[91][6] ),
    .S0(_06810_),
    .S1(_06811_),
    .X(_02692_));
 sky130_fd_sc_hd__o221a_1 _13611_ (.A1(_02689_),
    .A2(_02691_),
    .B1(_02692_),
    .B2(_06599_),
    .C1(_07219_),
    .X(_02693_));
 sky130_fd_sc_hd__mux4_1 _13612_ (.A0(\fifo0.fifo_store[80][6] ),
    .A1(\fifo0.fifo_store[81][6] ),
    .A2(\fifo0.fifo_store[82][6] ),
    .A3(\fifo0.fifo_store[83][6] ),
    .S0(_06450_),
    .S1(_06436_),
    .X(_02694_));
 sky130_fd_sc_hd__mux4_2 _13613_ (.A0(\fifo0.fifo_store[84][6] ),
    .A1(\fifo0.fifo_store[85][6] ),
    .A2(\fifo0.fifo_store[86][6] ),
    .A3(\fifo0.fifo_store[87][6] ),
    .S0(_06450_),
    .S1(_06436_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _13614_ (.A0(_02694_),
    .A1(_02695_),
    .S(_06440_),
    .X(_02696_));
 sky130_fd_sc_hd__a21o_1 _13615_ (.A1(_06868_),
    .A2(_02696_),
    .B1(_06493_),
    .X(_02697_));
 sky130_fd_sc_hd__mux4_1 _13616_ (.A0(\fifo0.fifo_store[76][6] ),
    .A1(\fifo0.fifo_store[77][6] ),
    .A2(\fifo0.fifo_store[78][6] ),
    .A3(\fifo0.fifo_store[79][6] ),
    .S0(_06625_),
    .S1(_06489_),
    .X(_02698_));
 sky130_fd_sc_hd__mux4_1 _13617_ (.A0(\fifo0.fifo_store[72][6] ),
    .A1(\fifo0.fifo_store[73][6] ),
    .A2(\fifo0.fifo_store[74][6] ),
    .A3(\fifo0.fifo_store[75][6] ),
    .S0(_06478_),
    .S1(_06627_),
    .X(_02699_));
 sky130_fd_sc_hd__or2_1 _13618_ (.A(_06484_),
    .B(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__o211a_1 _13619_ (.A1(_07371_),
    .A2(_02698_),
    .B1(_02700_),
    .C1(_06630_),
    .X(_02701_));
 sky130_fd_sc_hd__mux4_1 _13620_ (.A0(\fifo0.fifo_store[68][6] ),
    .A1(\fifo0.fifo_store[69][6] ),
    .A2(\fifo0.fifo_store[70][6] ),
    .A3(\fifo0.fifo_store[71][6] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02702_));
 sky130_fd_sc_hd__or2_1 _13621_ (.A(_06476_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__mux4_1 _13622_ (.A0(\fifo0.fifo_store[64][6] ),
    .A1(\fifo0.fifo_store[65][6] ),
    .A2(\fifo0.fifo_store[66][6] ),
    .A3(\fifo0.fifo_store[67][6] ),
    .S0(_06450_),
    .S1(_06436_),
    .X(_02704_));
 sky130_fd_sc_hd__or2_1 _13623_ (.A(_06447_),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__a31o_1 _13624_ (.A1(_06621_),
    .A2(_02703_),
    .A3(_02705_),
    .B1(_06641_),
    .X(_02706_));
 sky130_fd_sc_hd__o221a_1 _13625_ (.A1(_02693_),
    .A2(_02697_),
    .B1(_02701_),
    .B2(_02706_),
    .C1(_06497_),
    .X(_02707_));
 sky130_fd_sc_hd__a311o_4 _13626_ (.A1(_06465_),
    .A2(_02677_),
    .A3(_02687_),
    .B1(_02707_),
    .C1(_06604_),
    .X(_02708_));
 sky130_fd_sc_hd__mux4_1 _13627_ (.A0(\fifo0.fifo_store[0][6] ),
    .A1(\fifo0.fifo_store[1][6] ),
    .A2(\fifo0.fifo_store[2][6] ),
    .A3(\fifo0.fifo_store[3][6] ),
    .S0(_06479_),
    .S1(_06811_),
    .X(_02709_));
 sky130_fd_sc_hd__mux4_1 _13628_ (.A0(\fifo0.fifo_store[4][6] ),
    .A1(\fifo0.fifo_store[5][6] ),
    .A2(\fifo0.fifo_store[6][6] ),
    .A3(\fifo0.fifo_store[7][6] ),
    .S0(_06810_),
    .S1(_06811_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(_02709_),
    .A1(_02710_),
    .S(_06441_),
    .X(_02711_));
 sky130_fd_sc_hd__or2_1 _13630_ (.A(_06645_),
    .B(\fifo0.fifo_store[14][6] ),
    .X(_02712_));
 sky130_fd_sc_hd__o211a_1 _13631_ (.A1(_06612_),
    .A2(\fifo0.fifo_store[15][6] ),
    .B1(_02712_),
    .C1(_06648_),
    .X(_02713_));
 sky130_fd_sc_hd__mux2_1 _13632_ (.A0(\fifo0.fifo_store[12][6] ),
    .A1(\fifo0.fifo_store[13][6] ),
    .S(_06415_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_1 _13633_ (.A1(_06829_),
    .A2(_02714_),
    .B1(_06660_),
    .X(_02715_));
 sky130_fd_sc_hd__mux4_2 _13634_ (.A0(\fifo0.fifo_store[8][6] ),
    .A1(\fifo0.fifo_store[9][6] ),
    .A2(\fifo0.fifo_store[10][6] ),
    .A3(\fifo0.fifo_store[11][6] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_02716_));
 sky130_fd_sc_hd__o221a_1 _13635_ (.A1(_02713_),
    .A2(_02715_),
    .B1(_02716_),
    .B2(_06485_),
    .C1(_07219_),
    .X(_02717_));
 sky130_fd_sc_hd__a211o_1 _13636_ (.A1(_06793_),
    .A2(_02711_),
    .B1(_02717_),
    .C1(_06804_),
    .X(_02718_));
 sky130_fd_sc_hd__mux4_1 _13637_ (.A0(\fifo0.fifo_store[20][6] ),
    .A1(\fifo0.fifo_store[21][6] ),
    .A2(\fifo0.fifo_store[22][6] ),
    .A3(\fifo0.fifo_store[23][6] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_02719_));
 sky130_fd_sc_hd__or2_1 _13638_ (.A(_06456_),
    .B(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__mux4_1 _13639_ (.A0(\fifo0.fifo_store[16][6] ),
    .A1(\fifo0.fifo_store[17][6] ),
    .A2(\fifo0.fifo_store[18][6] ),
    .A3(\fifo0.fifo_store[19][6] ),
    .S0(_06533_),
    .S1(_06458_),
    .X(_02721_));
 sky130_fd_sc_hd__or2_1 _13640_ (.A(_06448_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__mux4_1 _13641_ (.A0(\fifo0.fifo_store[28][6] ),
    .A1(\fifo0.fifo_store[29][6] ),
    .A2(\fifo0.fifo_store[30][6] ),
    .A3(\fifo0.fifo_store[31][6] ),
    .S0(_07263_),
    .S1(_07391_),
    .X(_02723_));
 sky130_fd_sc_hd__mux4_1 _13642_ (.A0(\fifo0.fifo_store[24][6] ),
    .A1(\fifo0.fifo_store[25][6] ),
    .A2(\fifo0.fifo_store[26][6] ),
    .A3(\fifo0.fifo_store[27][6] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02724_));
 sky130_fd_sc_hd__or2_1 _13643_ (.A(_06447_),
    .B(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_1 _13644_ (.A1(_07371_),
    .A2(_02723_),
    .B1(_02725_),
    .C1(_07219_),
    .X(_02726_));
 sky130_fd_sc_hd__a311o_1 _13645_ (.A1(_06468_),
    .A2(_02720_),
    .A3(_02722_),
    .B1(_06539_),
    .C1(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__mux4_1 _13646_ (.A0(\fifo0.fifo_store[36][6] ),
    .A1(\fifo0.fifo_store[37][6] ),
    .A2(\fifo0.fifo_store[38][6] ),
    .A3(\fifo0.fifo_store[39][6] ),
    .S0(_07017_),
    .S1(_07391_),
    .X(_02728_));
 sky130_fd_sc_hd__mux4_1 _13647_ (.A0(\fifo0.fifo_store[32][6] ),
    .A1(\fifo0.fifo_store[33][6] ),
    .A2(\fifo0.fifo_store[34][6] ),
    .A3(\fifo0.fifo_store[35][6] ),
    .S0(_06520_),
    .S1(_06522_),
    .X(_02729_));
 sky130_fd_sc_hd__or2_1 _13648_ (.A(_06447_),
    .B(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__o211a_1 _13649_ (.A1(_07371_),
    .A2(_02728_),
    .B1(_02730_),
    .C1(_06868_),
    .X(_02731_));
 sky130_fd_sc_hd__mux4_1 _13650_ (.A0(\fifo0.fifo_store[40][6] ),
    .A1(\fifo0.fifo_store[41][6] ),
    .A2(\fifo0.fifo_store[42][6] ),
    .A3(\fifo0.fifo_store[43][6] ),
    .S0(_06848_),
    .S1(_06579_),
    .X(_02732_));
 sky130_fd_sc_hd__or2b_1 _13651_ (.A(\fifo0.fifo_store[47][6] ),
    .B_N(_06977_),
    .X(_02733_));
 sky130_fd_sc_hd__o21a_1 _13652_ (.A1(_06499_),
    .A2(\fifo0.fifo_store[46][6] ),
    .B1(_06647_),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _13653_ (.A0(\fifo0.fifo_store[44][6] ),
    .A1(\fifo0.fifo_store[45][6] ),
    .S(_06415_),
    .X(_02735_));
 sky130_fd_sc_hd__a221o_1 _13654_ (.A1(_02733_),
    .A2(_02734_),
    .B1(_02735_),
    .B2(_06650_),
    .C1(_06660_),
    .X(_02736_));
 sky130_fd_sc_hd__o211a_1 _13655_ (.A1(_06624_),
    .A2(_02732_),
    .B1(_02736_),
    .C1(_06630_),
    .X(_02737_));
 sky130_fd_sc_hd__mux4_2 _13656_ (.A0(\fifo0.fifo_store[52][6] ),
    .A1(\fifo0.fifo_store[53][6] ),
    .A2(\fifo0.fifo_store[54][6] ),
    .A3(\fifo0.fifo_store[55][6] ),
    .S0(_06450_),
    .S1(_06436_),
    .X(_02738_));
 sky130_fd_sc_hd__mux4_1 _13657_ (.A0(\fifo0.fifo_store[48][6] ),
    .A1(\fifo0.fifo_store[49][6] ),
    .A2(\fifo0.fifo_store[50][6] ),
    .A3(\fifo0.fifo_store[51][6] ),
    .S0(_06450_),
    .S1(_06436_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(_02738_),
    .A1(_02739_),
    .S(_06430_),
    .X(_02740_));
 sky130_fd_sc_hd__mux4_1 _13659_ (.A0(\fifo0.fifo_store[56][6] ),
    .A1(\fifo0.fifo_store[57][6] ),
    .A2(\fifo0.fifo_store[58][6] ),
    .A3(\fifo0.fifo_store[59][6] ),
    .S0(_06426_),
    .S1(_06488_),
    .X(_02741_));
 sky130_fd_sc_hd__or2_1 _13660_ (.A(_06623_),
    .B(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__mux4_2 _13661_ (.A0(\fifo0.fifo_store[60][6] ),
    .A1(\fifo0.fifo_store[61][6] ),
    .A2(\fifo0.fifo_store[62][6] ),
    .A3(\fifo0.fifo_store[63][6] ),
    .S0(_06657_),
    .S1(_06510_),
    .X(_02743_));
 sky130_fd_sc_hd__o21a_1 _13662_ (.A1(_06668_),
    .A2(_02743_),
    .B1(_06461_),
    .X(_02744_));
 sky130_fd_sc_hd__a221o_1 _13663_ (.A1(_06868_),
    .A2(_02740_),
    .B1(_02742_),
    .B2(_02744_),
    .C1(_06493_),
    .X(_02745_));
 sky130_fd_sc_hd__o311a_1 _13664_ (.A1(_06589_),
    .A2(_02731_),
    .A3(_02737_),
    .B1(_02745_),
    .C1(_06643_),
    .X(_02746_));
 sky130_fd_sc_hd__a311o_2 _13665_ (.A1(_06575_),
    .A2(_02718_),
    .A3(_02727_),
    .B1(_00006_),
    .C1(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__nor2_1 _13666_ (.A(_06391_),
    .B(_06774_),
    .Y(_02748_));
 sky130_fd_sc_hd__o221a_1 _13667_ (.A1(_06396_),
    .A2(_02748_),
    .B1(_06920_),
    .B2(_06912_),
    .C1(_06358_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _13668_ (.A(_02165_),
    .B(_06784_),
    .X(_02750_));
 sky130_fd_sc_hd__o21a_1 _13669_ (.A1(_06888_),
    .A2(_02750_),
    .B1(_06401_),
    .X(_02751_));
 sky130_fd_sc_hd__o21a_1 _13670_ (.A1(_02749_),
    .A2(_02751_),
    .B1(_06747_),
    .X(_02752_));
 sky130_fd_sc_hd__a21oi_1 _13671_ (.A1(_06378_),
    .A2(_06779_),
    .B1(_06760_),
    .Y(_02753_));
 sky130_fd_sc_hd__nor3_1 _13672_ (.A(_06747_),
    .B(_02749_),
    .C(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__or2_1 _13673_ (.A(\sinegen0.read_ptr[4] ),
    .B(_06891_),
    .X(_02755_));
 sky130_fd_sc_hd__a21o_1 _13674_ (.A1(_06377_),
    .A2(_06786_),
    .B1(_06923_),
    .X(_02756_));
 sky130_fd_sc_hd__o21a_1 _13675_ (.A1(_06393_),
    .A2(_07056_),
    .B1(\sinegen0.read_ptr[4] ),
    .X(_02757_));
 sky130_fd_sc_hd__a2bb2o_1 _13676_ (.A1_N(_07431_),
    .A2_N(_02755_),
    .B1(_02756_),
    .B2(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__a31o_1 _13677_ (.A1(_06363_),
    .A2(_06384_),
    .A3(_06766_),
    .B1(_02755_),
    .X(_02759_));
 sky130_fd_sc_hd__a21oi_1 _13678_ (.A1(_02756_),
    .A2(_02757_),
    .B1(\sinegen0.read_ptr[6] ),
    .Y(_02760_));
 sky130_fd_sc_hd__a221o_1 _13679_ (.A1(\sinegen0.read_ptr[6] ),
    .A2(_02758_),
    .B1(_02759_),
    .B2(_02760_),
    .C1(_06370_),
    .X(_02761_));
 sky130_fd_sc_hd__o311a_1 _13680_ (.A1(_06405_),
    .A2(_02752_),
    .A3(_02754_),
    .B1(net23),
    .C1(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__a31o_1 _13681_ (.A1(_06606_),
    .A2(_02708_),
    .A3(_02747_),
    .B1(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _13682_ (.A0(_02668_),
    .A1(_02763_),
    .S(_06353_),
    .X(_02764_));
 sky130_fd_sc_hd__mux4_1 _13683_ (.A0(_02177_),
    .A1(_02179_),
    .A2(_02574_),
    .A3(_02764_),
    .S0(_07315_),
    .S1(_07326_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _13684_ (.A0(_02385_),
    .A1(_02765_),
    .S(_07314_),
    .X(_02766_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(_02383_),
    .B(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__and2_1 _13686_ (.A(_02382_),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__nor2_1 _13687_ (.A(_02382_),
    .B(_02767_),
    .Y(_02769_));
 sky130_fd_sc_hd__or2_1 _13688_ (.A(_02768_),
    .B(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _13689_ (.A0(_02174_),
    .A1(_02177_),
    .S(_07315_),
    .X(_02771_));
 sky130_fd_sc_hd__mux2_1 _13690_ (.A0(_02179_),
    .A1(_02574_),
    .S(_07315_),
    .X(_02772_));
 sky130_fd_sc_hd__mux4_2 _13691_ (.A0(\fifo0.fifo_store[60][4] ),
    .A1(\fifo0.fifo_store[61][4] ),
    .A2(\fifo0.fifo_store[62][4] ),
    .A3(\fifo0.fifo_store[63][4] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_02773_));
 sky130_fd_sc_hd__mux4_1 _13692_ (.A0(\fifo0.fifo_store[56][4] ),
    .A1(\fifo0.fifo_store[57][4] ),
    .A2(\fifo0.fifo_store[58][4] ),
    .A3(\fifo0.fifo_store[59][4] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_02774_));
 sky130_fd_sc_hd__or2_1 _13693_ (.A(_06797_),
    .B(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__o211a_1 _13694_ (.A1(_07355_),
    .A2(_02773_),
    .B1(_02775_),
    .C1(_07094_),
    .X(_02776_));
 sky130_fd_sc_hd__mux4_1 _13695_ (.A0(\fifo0.fifo_store[48][4] ),
    .A1(\fifo0.fifo_store[49][4] ),
    .A2(\fifo0.fifo_store[50][4] ),
    .A3(\fifo0.fifo_store[51][4] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_02777_));
 sky130_fd_sc_hd__or2b_1 _13696_ (.A(\fifo0.fifo_store[55][4] ),
    .B_N(_07067_),
    .X(_02778_));
 sky130_fd_sc_hd__o21a_1 _13697_ (.A1(_07067_),
    .A2(\fifo0.fifo_store[54][4] ),
    .B1(_06481_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(\fifo0.fifo_store[52][4] ),
    .A1(\fifo0.fifo_store[53][4] ),
    .S(_06870_),
    .X(_02780_));
 sky130_fd_sc_hd__a221o_1 _13699_ (.A1(_02778_),
    .A2(_02779_),
    .B1(_02780_),
    .B2(_06516_),
    .C1(_07132_),
    .X(_02781_));
 sky130_fd_sc_hd__o211a_1 _13700_ (.A1(_06442_),
    .A2(_02777_),
    .B1(_02781_),
    .C1(_06552_),
    .X(_02782_));
 sky130_fd_sc_hd__mux4_1 _13701_ (.A0(\fifo0.fifo_store[40][4] ),
    .A1(\fifo0.fifo_store[41][4] ),
    .A2(\fifo0.fifo_store[42][4] ),
    .A3(\fifo0.fifo_store[43][4] ),
    .S0(_06977_),
    .S1(_06437_),
    .X(_02783_));
 sky130_fd_sc_hd__or2_1 _13702_ (.A(_06441_),
    .B(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__mux4_2 _13703_ (.A0(\fifo0.fifo_store[44][4] ),
    .A1(\fifo0.fifo_store[45][4] ),
    .A2(\fifo0.fifo_store[46][4] ),
    .A3(\fifo0.fifo_store[47][4] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_02785_));
 sky130_fd_sc_hd__o21a_1 _13704_ (.A1(_06502_),
    .A2(_02785_),
    .B1(_06462_),
    .X(_02786_));
 sky130_fd_sc_hd__mux4_1 _13705_ (.A0(\fifo0.fifo_store[36][4] ),
    .A1(\fifo0.fifo_store[37][4] ),
    .A2(\fifo0.fifo_store[38][4] ),
    .A3(\fifo0.fifo_store[39][4] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_02787_));
 sky130_fd_sc_hd__or2_1 _13706_ (.A(_06456_),
    .B(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__mux4_1 _13707_ (.A0(\fifo0.fifo_store[32][4] ),
    .A1(\fifo0.fifo_store[33][4] ),
    .A2(\fifo0.fifo_store[34][4] ),
    .A3(\fifo0.fifo_store[35][4] ),
    .S0(_06521_),
    .S1(_06555_),
    .X(_02789_));
 sky130_fd_sc_hd__o21a_1 _13708_ (.A1(_06519_),
    .A2(_02789_),
    .B1(_06467_),
    .X(_02790_));
 sky130_fd_sc_hd__a221o_1 _13709_ (.A1(_02784_),
    .A2(_02786_),
    .B1(_02788_),
    .B2(_02790_),
    .C1(_06408_),
    .X(_02791_));
 sky130_fd_sc_hd__o311a_1 _13710_ (.A1(_07085_),
    .A2(_02776_),
    .A3(_02782_),
    .B1(_06465_),
    .C1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__or2_1 _13711_ (.A(_07001_),
    .B(\fifo0.fifo_store[6][4] ),
    .X(_02793_));
 sky130_fd_sc_hd__o211a_1 _13712_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[7][4] ),
    .B1(_02793_),
    .C1(_07257_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _13713_ (.A0(\fifo0.fifo_store[4][4] ),
    .A1(\fifo0.fifo_store[5][4] ),
    .S(_06870_),
    .X(_02795_));
 sky130_fd_sc_hd__a21o_1 _13714_ (.A1(_06516_),
    .A2(_02795_),
    .B1(_07132_),
    .X(_02796_));
 sky130_fd_sc_hd__mux4_1 _13715_ (.A0(\fifo0.fifo_store[0][4] ),
    .A1(\fifo0.fifo_store[1][4] ),
    .A2(\fifo0.fifo_store[2][4] ),
    .A3(\fifo0.fifo_store[3][4] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_02797_));
 sky130_fd_sc_hd__o221a_1 _13716_ (.A1(_02794_),
    .A2(_02796_),
    .B1(_02797_),
    .B2(_06442_),
    .C1(_06445_),
    .X(_02798_));
 sky130_fd_sc_hd__mux4_2 _13717_ (.A0(\fifo0.fifo_store[8][4] ),
    .A1(\fifo0.fifo_store[9][4] ),
    .A2(\fifo0.fifo_store[10][4] ),
    .A3(\fifo0.fifo_store[11][4] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_02799_));
 sky130_fd_sc_hd__mux4_1 _13718_ (.A0(\fifo0.fifo_store[12][4] ),
    .A1(\fifo0.fifo_store[13][4] ),
    .A2(\fifo0.fifo_store[14][4] ),
    .A3(\fifo0.fifo_store[15][4] ),
    .S0(_06499_),
    .S1(_06437_),
    .X(_02800_));
 sky130_fd_sc_hd__or2_1 _13719_ (.A(_06517_),
    .B(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__o211a_1 _13720_ (.A1(_06449_),
    .A2(_02799_),
    .B1(_02801_),
    .C1(_06463_),
    .X(_02802_));
 sky130_fd_sc_hd__mux4_1 _13721_ (.A0(\fifo0.fifo_store[16][4] ),
    .A1(\fifo0.fifo_store[17][4] ),
    .A2(\fifo0.fifo_store[18][4] ),
    .A3(\fifo0.fifo_store[19][4] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_02803_));
 sky130_fd_sc_hd__mux4_1 _13722_ (.A0(\fifo0.fifo_store[20][4] ),
    .A1(\fifo0.fifo_store[21][4] ),
    .A2(\fifo0.fifo_store[22][4] ),
    .A3(\fifo0.fifo_store[23][4] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _13723_ (.A0(_02803_),
    .A1(_02804_),
    .S(_06565_),
    .X(_02805_));
 sky130_fd_sc_hd__mux4_1 _13724_ (.A0(\fifo0.fifo_store[28][4] ),
    .A1(\fifo0.fifo_store[29][4] ),
    .A2(\fifo0.fifo_store[30][4] ),
    .A3(\fifo0.fifo_store[31][4] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_02806_));
 sky130_fd_sc_hd__or2_1 _13725_ (.A(_06456_),
    .B(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__mux4_1 _13726_ (.A0(\fifo0.fifo_store[24][4] ),
    .A1(\fifo0.fifo_store[25][4] ),
    .A2(\fifo0.fifo_store[26][4] ),
    .A3(\fifo0.fifo_store[27][4] ),
    .S0(_06521_),
    .S1(_06555_),
    .X(_02808_));
 sky130_fd_sc_hd__o21a_1 _13727_ (.A1(_06599_),
    .A2(_02808_),
    .B1(_06571_),
    .X(_02809_));
 sky130_fd_sc_hd__a221o_1 _13728_ (.A1(_06552_),
    .A2(_02805_),
    .B1(_02807_),
    .B2(_02809_),
    .C1(_06539_),
    .X(_02810_));
 sky130_fd_sc_hd__o311a_1 _13729_ (.A1(_06409_),
    .A2(_02798_),
    .A3(_02802_),
    .B1(_02810_),
    .C1(_06498_),
    .X(_02811_));
 sky130_fd_sc_hd__mux4_1 _13730_ (.A0(\fifo0.fifo_store[88][4] ),
    .A1(\fifo0.fifo_store[89][4] ),
    .A2(\fifo0.fifo_store[90][4] ),
    .A3(\fifo0.fifo_store[91][4] ),
    .S0(_06536_),
    .S1(_06523_),
    .X(_02812_));
 sky130_fd_sc_hd__or2_1 _13731_ (.A(_06519_),
    .B(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__mux4_2 _13732_ (.A0(\fifo0.fifo_store[92][4] ),
    .A1(\fifo0.fifo_store[93][4] ),
    .A2(\fifo0.fifo_store[94][4] ),
    .A3(\fifo0.fifo_store[95][4] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_02814_));
 sky130_fd_sc_hd__o21a_1 _13733_ (.A1(_06477_),
    .A2(_02814_),
    .B1(_06571_),
    .X(_02815_));
 sky130_fd_sc_hd__mux4_1 _13734_ (.A0(\fifo0.fifo_store[84][4] ),
    .A1(\fifo0.fifo_store[85][4] ),
    .A2(\fifo0.fifo_store[86][4] ),
    .A3(\fifo0.fifo_store[87][4] ),
    .S0(_06810_),
    .S1(_06555_),
    .X(_02816_));
 sky130_fd_sc_hd__or2_1 _13735_ (.A(_06477_),
    .B(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__mux4_1 _13736_ (.A0(\fifo0.fifo_store[80][4] ),
    .A1(\fifo0.fifo_store[81][4] ),
    .A2(\fifo0.fifo_store[82][4] ),
    .A3(\fifo0.fifo_store[83][4] ),
    .S0(_07017_),
    .S1(_07391_),
    .X(_02818_));
 sky130_fd_sc_hd__o21a_1 _13737_ (.A1(_06485_),
    .A2(_02818_),
    .B1(_06467_),
    .X(_02819_));
 sky130_fd_sc_hd__a221o_1 _13738_ (.A1(_02813_),
    .A2(_02815_),
    .B1(_02817_),
    .B2(_02819_),
    .C1(_06494_),
    .X(_02820_));
 sky130_fd_sc_hd__or2b_1 _13739_ (.A(\fifo0.fifo_store[79][4] ),
    .B_N(_07097_),
    .X(_02821_));
 sky130_fd_sc_hd__o21a_1 _13740_ (.A1(_07097_),
    .A2(\fifo0.fifo_store[78][4] ),
    .B1(_06421_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _13741_ (.A0(\fifo0.fifo_store[76][4] ),
    .A1(\fifo0.fifo_store[77][4] ),
    .S(_06946_),
    .X(_02823_));
 sky130_fd_sc_hd__a221o_1 _13742_ (.A1(_02821_),
    .A2(_02822_),
    .B1(_02823_),
    .B2(_06425_),
    .C1(_06477_),
    .X(_02824_));
 sky130_fd_sc_hd__mux4_1 _13743_ (.A0(\fifo0.fifo_store[72][4] ),
    .A1(\fifo0.fifo_store[73][4] ),
    .A2(\fifo0.fifo_store[74][4] ),
    .A3(\fifo0.fifo_store[75][4] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_02825_));
 sky130_fd_sc_hd__o21a_1 _13744_ (.A1(_06485_),
    .A2(_02825_),
    .B1(_06571_),
    .X(_02826_));
 sky130_fd_sc_hd__mux4_2 _13745_ (.A0(\fifo0.fifo_store[64][4] ),
    .A1(\fifo0.fifo_store[65][4] ),
    .A2(\fifo0.fifo_store[66][4] ),
    .A3(\fifo0.fifo_store[67][4] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_02827_));
 sky130_fd_sc_hd__mux4_1 _13746_ (.A0(\fifo0.fifo_store[68][4] ),
    .A1(\fifo0.fifo_store[69][4] ),
    .A2(\fifo0.fifo_store[70][4] ),
    .A3(\fifo0.fifo_store[71][4] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(_02827_),
    .A1(_02828_),
    .S(_06797_),
    .X(_02829_));
 sky130_fd_sc_hd__a221o_1 _13748_ (.A1(_02824_),
    .A2(_02826_),
    .B1(_02829_),
    .B2(_06468_),
    .C1(_06589_),
    .X(_02830_));
 sky130_fd_sc_hd__and3_1 _13749_ (.A(_06575_),
    .B(_02820_),
    .C(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__or2b_1 _13750_ (.A(\fifo0.fifo_store[127][4] ),
    .B_N(_06542_),
    .X(_02832_));
 sky130_fd_sc_hd__o21a_1 _13751_ (.A1(_06435_),
    .A2(\fifo0.fifo_store[126][4] ),
    .B1(_06615_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _13752_ (.A0(\fifo0.fifo_store[124][4] ),
    .A1(\fifo0.fifo_store[125][4] ),
    .S(_07001_),
    .X(_02834_));
 sky130_fd_sc_hd__a221o_1 _13753_ (.A1(_02832_),
    .A2(_02833_),
    .B1(_02834_),
    .B2(_06954_),
    .C1(_06477_),
    .X(_02835_));
 sky130_fd_sc_hd__mux4_2 _13754_ (.A0(\fifo0.fifo_store[120][4] ),
    .A1(\fifo0.fifo_store[121][4] ),
    .A2(\fifo0.fifo_store[122][4] ),
    .A3(\fifo0.fifo_store[123][4] ),
    .S0(_06693_),
    .S1(_06579_),
    .X(_02836_));
 sky130_fd_sc_hd__o21a_1 _13755_ (.A1(_06624_),
    .A2(_02836_),
    .B1(_07219_),
    .X(_02837_));
 sky130_fd_sc_hd__mux4_1 _13756_ (.A0(\fifo0.fifo_store[112][4] ),
    .A1(\fifo0.fifo_store[113][4] ),
    .A2(\fifo0.fifo_store[114][4] ),
    .A3(\fifo0.fifo_store[115][4] ),
    .S0(_06600_),
    .S1(_06555_),
    .X(_02838_));
 sky130_fd_sc_hd__mux4_1 _13757_ (.A0(\fifo0.fifo_store[116][4] ),
    .A1(\fifo0.fifo_store[117][4] ),
    .A2(\fifo0.fifo_store[118][4] ),
    .A3(\fifo0.fifo_store[119][4] ),
    .S0(_06600_),
    .S1(_06555_),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _13758_ (.A0(_02838_),
    .A1(_02839_),
    .S(_06441_),
    .X(_02840_));
 sky130_fd_sc_hd__a221o_1 _13759_ (.A1(_02835_),
    .A2(_02837_),
    .B1(_02840_),
    .B2(_06793_),
    .C1(_06494_),
    .X(_02841_));
 sky130_fd_sc_hd__mux4_2 _13760_ (.A0(\fifo0.fifo_store[104][4] ),
    .A1(\fifo0.fifo_store[105][4] ),
    .A2(\fifo0.fifo_store[106][4] ),
    .A3(\fifo0.fifo_store[107][4] ),
    .S0(_07263_),
    .S1(_06481_),
    .X(_02842_));
 sky130_fd_sc_hd__or2_1 _13761_ (.A(_06599_),
    .B(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__mux4_1 _13762_ (.A0(\fifo0.fifo_store[108][4] ),
    .A1(\fifo0.fifo_store[109][4] ),
    .A2(\fifo0.fifo_store[110][4] ),
    .A3(\fifo0.fifo_store[111][4] ),
    .S0(_06625_),
    .S1(_06489_),
    .X(_02844_));
 sky130_fd_sc_hd__o21a_1 _13763_ (.A1(_07371_),
    .A2(_02844_),
    .B1(_07219_),
    .X(_02845_));
 sky130_fd_sc_hd__mux4_2 _13764_ (.A0(\fifo0.fifo_store[96][4] ),
    .A1(\fifo0.fifo_store[97][4] ),
    .A2(\fifo0.fifo_store[98][4] ),
    .A3(\fifo0.fifo_store[99][4] ),
    .S0(_06487_),
    .S1(_07391_),
    .X(_02846_));
 sky130_fd_sc_hd__or2_1 _13765_ (.A(_06485_),
    .B(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__mux4_1 _13766_ (.A0(\fifo0.fifo_store[100][4] ),
    .A1(\fifo0.fifo_store[101][4] ),
    .A2(\fifo0.fifo_store[102][4] ),
    .A3(\fifo0.fifo_store[103][4] ),
    .S0(_06658_),
    .S1(_06511_),
    .X(_02848_));
 sky130_fd_sc_hd__o21a_1 _13767_ (.A1(_06814_),
    .A2(_02848_),
    .B1(_06868_),
    .X(_02849_));
 sky130_fd_sc_hd__a221o_1 _13768_ (.A1(_02843_),
    .A2(_02845_),
    .B1(_02847_),
    .B2(_02849_),
    .C1(_06804_),
    .X(_02850_));
 sky130_fd_sc_hd__a31o_1 _13769_ (.A1(_06792_),
    .A2(_02841_),
    .A3(_02850_),
    .B1(_06604_),
    .X(_02851_));
 sky130_fd_sc_hd__o32a_2 _13770_ (.A1(_06992_),
    .A2(_02792_),
    .A3(_02811_),
    .B1(_02831_),
    .B2(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a21o_1 _13771_ (.A1(_06764_),
    .A2(_06781_),
    .B1(_06922_),
    .X(_02853_));
 sky130_fd_sc_hd__a21oi_1 _13772_ (.A1(_06768_),
    .A2(_02853_),
    .B1(_07198_),
    .Y(_02854_));
 sky130_fd_sc_hd__nand2_1 _13773_ (.A(_06922_),
    .B(_06781_),
    .Y(_02855_));
 sky130_fd_sc_hd__or2b_1 _13774_ (.A(_06373_),
    .B_N(_06404_),
    .X(_02856_));
 sky130_fd_sc_hd__nor4_1 _13775_ (.A(_06392_),
    .B(_06387_),
    .C(_02856_),
    .D(_06393_),
    .Y(_02857_));
 sky130_fd_sc_hd__and3b_1 _13776_ (.A_N(_06392_),
    .B(_02165_),
    .C(_06910_),
    .X(_02858_));
 sky130_fd_sc_hd__a311o_1 _13777_ (.A1(_07193_),
    .A2(_02853_),
    .A3(_02855_),
    .B1(_02857_),
    .C1(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__o21ai_1 _13778_ (.A1(_02854_),
    .A2(_02859_),
    .B1(_06769_),
    .Y(_02860_));
 sky130_fd_sc_hd__o311a_1 _13779_ (.A1(_02666_),
    .A2(_02854_),
    .A3(_02859_),
    .B1(_02860_),
    .C1(_06918_),
    .X(_02861_));
 sky130_fd_sc_hd__a211o_1 _13780_ (.A1(_06611_),
    .A2(_02852_),
    .B1(_02861_),
    .C1(_07163_),
    .X(_02862_));
 sky130_fd_sc_hd__buf_8 _13781_ (.A(_06542_),
    .X(_02863_));
 sky130_fd_sc_hd__buf_6 _13782_ (.A(_07099_),
    .X(_02864_));
 sky130_fd_sc_hd__mux4_1 _13783_ (.A0(\fifo0.fifo_store[72][3] ),
    .A1(\fifo0.fifo_store[73][3] ),
    .A2(\fifo0.fifo_store[74][3] ),
    .A3(\fifo0.fifo_store[75][3] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__buf_4 _13784_ (.A(_07371_),
    .X(_02866_));
 sky130_fd_sc_hd__buf_8 _13785_ (.A(_06693_),
    .X(_02867_));
 sky130_fd_sc_hd__mux4_1 _13786_ (.A0(\fifo0.fifo_store[76][3] ),
    .A1(\fifo0.fifo_store[77][3] ),
    .A2(\fifo0.fifo_store[78][3] ),
    .A3(\fifo0.fifo_store[79][3] ),
    .S0(_02867_),
    .S1(_07257_),
    .X(_02868_));
 sky130_fd_sc_hd__o21a_1 _13787_ (.A1(_02866_),
    .A2(_02868_),
    .B1(_06463_),
    .X(_02869_));
 sky130_fd_sc_hd__o21ai_2 _13788_ (.A1(_07203_),
    .A2(_02865_),
    .B1(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__buf_8 _13789_ (.A(_07022_),
    .X(_02871_));
 sky130_fd_sc_hd__or2_1 _13790_ (.A(_02871_),
    .B(\fifo0.fifo_store[68][3] ),
    .X(_02872_));
 sky130_fd_sc_hd__o211a_1 _13791_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[69][3] ),
    .B1(_02872_),
    .C1(_06954_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _13792_ (.A0(\fifo0.fifo_store[70][3] ),
    .A1(\fifo0.fifo_store[71][3] ),
    .S(_07079_),
    .X(_02874_));
 sky130_fd_sc_hd__a21o_1 _13793_ (.A1(_02864_),
    .A2(_02874_),
    .B1(_07355_),
    .X(_02875_));
 sky130_fd_sc_hd__mux4_2 _13794_ (.A0(\fifo0.fifo_store[64][3] ),
    .A1(\fifo0.fifo_store[65][3] ),
    .A2(\fifo0.fifo_store[66][3] ),
    .A3(\fifo0.fifo_store[67][3] ),
    .S0(_07204_),
    .S1(_02864_),
    .X(_02876_));
 sky130_fd_sc_hd__o221ai_1 _13795_ (.A1(_02873_),
    .A2(_02875_),
    .B1(_02876_),
    .B2(_07203_),
    .C1(_06939_),
    .Y(_02877_));
 sky130_fd_sc_hd__clkbuf_16 _13796_ (.A(_06569_),
    .X(_02878_));
 sky130_fd_sc_hd__buf_8 _13797_ (.A(_07391_),
    .X(_02879_));
 sky130_fd_sc_hd__mux4_1 _13798_ (.A0(\fifo0.fifo_store[88][3] ),
    .A1(\fifo0.fifo_store[89][3] ),
    .A2(\fifo0.fifo_store[90][3] ),
    .A3(\fifo0.fifo_store[91][3] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_06554_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__mux4_1 _13800_ (.A0(\fifo0.fifo_store[92][3] ),
    .A1(\fifo0.fifo_store[93][3] ),
    .A2(\fifo0.fifo_store[94][3] ),
    .A3(\fifo0.fifo_store[95][3] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_02882_));
 sky130_fd_sc_hd__o21ai_1 _13801_ (.A1(_07355_),
    .A2(_02882_),
    .B1(_06463_),
    .Y(_02883_));
 sky130_fd_sc_hd__mux4_1 _13802_ (.A0(\fifo0.fifo_store[84][3] ),
    .A1(\fifo0.fifo_store[85][3] ),
    .A2(\fifo0.fifo_store[86][3] ),
    .A3(\fifo0.fifo_store[87][3] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_02884_));
 sky130_fd_sc_hd__nor2_1 _13803_ (.A(_02866_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__mux4_1 _13804_ (.A0(\fifo0.fifo_store[80][3] ),
    .A1(\fifo0.fifo_store[81][3] ),
    .A2(\fifo0.fifo_store[82][3] ),
    .A3(\fifo0.fifo_store[83][3] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_02886_));
 sky130_fd_sc_hd__o21ai_1 _13805_ (.A1(_06449_),
    .A2(_02886_),
    .B1(_06468_),
    .Y(_02887_));
 sky130_fd_sc_hd__o221a_1 _13806_ (.A1(_02881_),
    .A2(_02883_),
    .B1(_02885_),
    .B2(_02887_),
    .C1(_06966_),
    .X(_02888_));
 sky130_fd_sc_hd__a311o_1 _13807_ (.A1(_07354_),
    .A2(_02870_),
    .A3(_02877_),
    .B1(_06792_),
    .C1(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__mux4_2 _13808_ (.A0(\fifo0.fifo_store[120][3] ),
    .A1(\fifo0.fifo_store[121][3] ),
    .A2(\fifo0.fifo_store[122][3] ),
    .A3(\fifo0.fifo_store[123][3] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_02890_));
 sky130_fd_sc_hd__mux4_1 _13809_ (.A0(\fifo0.fifo_store[124][3] ),
    .A1(\fifo0.fifo_store[125][3] ),
    .A2(\fifo0.fifo_store[126][3] ),
    .A3(\fifo0.fifo_store[127][3] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_02891_));
 sky130_fd_sc_hd__o21a_1 _13810_ (.A1(_02866_),
    .A2(_02891_),
    .B1(_07220_),
    .X(_02892_));
 sky130_fd_sc_hd__o21ai_1 _13811_ (.A1(_07203_),
    .A2(_02890_),
    .B1(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__buf_4 _13812_ (.A(_06797_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _13813_ (.A0(\fifo0.fifo_store[116][3] ),
    .A1(\fifo0.fifo_store[117][3] ),
    .S(_02871_),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_1 _13814_ (.A(_07207_),
    .B(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__buf_4 _13815_ (.A(_07205_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _13816_ (.A0(\fifo0.fifo_store[118][3] ),
    .A1(\fifo0.fifo_store[119][3] ),
    .S(_02871_),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _13817_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__mux4_1 _13818_ (.A0(\fifo0.fifo_store[112][3] ),
    .A1(\fifo0.fifo_store[113][3] ),
    .A2(\fifo0.fifo_store[114][3] ),
    .A3(\fifo0.fifo_store[115][3] ),
    .S0(_06452_),
    .S1(_06556_),
    .X(_02900_));
 sky130_fd_sc_hd__o21ai_1 _13819_ (.A1(_06449_),
    .A2(_02900_),
    .B1(_06468_),
    .Y(_02901_));
 sky130_fd_sc_hd__a31o_1 _13820_ (.A1(_02894_),
    .A2(_02896_),
    .A3(_02899_),
    .B1(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__mux4_1 _13821_ (.A0(\fifo0.fifo_store[104][3] ),
    .A1(\fifo0.fifo_store[105][3] ),
    .A2(\fifo0.fifo_store[106][3] ),
    .A3(\fifo0.fifo_store[107][3] ),
    .S0(_06951_),
    .S1(_06556_),
    .X(_02903_));
 sky130_fd_sc_hd__nor2_1 _13822_ (.A(_06449_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__mux4_1 _13823_ (.A0(\fifo0.fifo_store[108][3] ),
    .A1(\fifo0.fifo_store[109][3] ),
    .A2(\fifo0.fifo_store[110][3] ),
    .A3(\fifo0.fifo_store[111][3] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_02905_));
 sky130_fd_sc_hd__o21ai_1 _13824_ (.A1(_07355_),
    .A2(_02905_),
    .B1(_07094_),
    .Y(_02906_));
 sky130_fd_sc_hd__mux4_2 _13825_ (.A0(\fifo0.fifo_store[100][3] ),
    .A1(\fifo0.fifo_store[101][3] ),
    .A2(\fifo0.fifo_store[102][3] ),
    .A3(\fifo0.fifo_store[103][3] ),
    .S0(_06951_),
    .S1(_02879_),
    .X(_02907_));
 sky130_fd_sc_hd__nor2_1 _13826_ (.A(_07355_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__mux4_1 _13827_ (.A0(\fifo0.fifo_store[96][3] ),
    .A1(\fifo0.fifo_store[97][3] ),
    .A2(\fifo0.fifo_store[98][3] ),
    .A3(\fifo0.fifo_store[99][3] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_02909_));
 sky130_fd_sc_hd__o21ai_2 _13828_ (.A1(_06442_),
    .A2(_02909_),
    .B1(_06552_),
    .Y(_02910_));
 sky130_fd_sc_hd__o221a_1 _13829_ (.A1(_02904_),
    .A2(_02906_),
    .B1(_02908_),
    .B2(_02910_),
    .C1(_07085_),
    .X(_02911_));
 sky130_fd_sc_hd__a311o_1 _13830_ (.A1(_07202_),
    .A2(_02893_),
    .A3(_02902_),
    .B1(_02911_),
    .C1(_06575_),
    .X(_02912_));
 sky130_fd_sc_hd__nand3_4 _13831_ (.A(_06992_),
    .B(_02889_),
    .C(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__or2_1 _13832_ (.A(_07001_),
    .B(\fifo0.fifo_store[6][3] ),
    .X(_02914_));
 sky130_fd_sc_hd__o211a_1 _13833_ (.A1(_06413_),
    .A2(\fifo0.fifo_store[7][3] ),
    .B1(_02914_),
    .C1(_07257_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _13834_ (.A0(\fifo0.fifo_store[4][3] ),
    .A1(\fifo0.fifo_store[5][3] ),
    .S(_06549_),
    .X(_02916_));
 sky130_fd_sc_hd__a21o_1 _13835_ (.A1(_06425_),
    .A2(_02916_),
    .B1(_06431_),
    .X(_02917_));
 sky130_fd_sc_hd__mux4_1 _13836_ (.A0(\fifo0.fifo_store[0][3] ),
    .A1(\fifo0.fifo_store[1][3] ),
    .A2(\fifo0.fifo_store[2][3] ),
    .A3(\fifo0.fifo_store[3][3] ),
    .S0(_06435_),
    .S1(_07099_),
    .X(_02918_));
 sky130_fd_sc_hd__o221a_1 _13837_ (.A1(_02915_),
    .A2(_02917_),
    .B1(_02918_),
    .B2(_06442_),
    .C1(_06445_),
    .X(_02919_));
 sky130_fd_sc_hd__mux4_2 _13838_ (.A0(\fifo0.fifo_store[8][3] ),
    .A1(\fifo0.fifo_store[9][3] ),
    .A2(\fifo0.fifo_store[10][3] ),
    .A3(\fifo0.fifo_store[11][3] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_02920_));
 sky130_fd_sc_hd__mux4_1 _13839_ (.A0(\fifo0.fifo_store[12][3] ),
    .A1(\fifo0.fifo_store[13][3] ),
    .A2(\fifo0.fifo_store[14][3] ),
    .A3(\fifo0.fifo_store[15][3] ),
    .S0(_06591_),
    .S1(_06592_),
    .X(_02921_));
 sky130_fd_sc_hd__or2_1 _13840_ (.A(_06517_),
    .B(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__o211a_1 _13841_ (.A1(_06449_),
    .A2(_02920_),
    .B1(_02922_),
    .C1(_06463_),
    .X(_02923_));
 sky130_fd_sc_hd__mux4_1 _13842_ (.A0(\fifo0.fifo_store[16][3] ),
    .A1(\fifo0.fifo_store[17][3] ),
    .A2(\fifo0.fifo_store[18][3] ),
    .A3(\fifo0.fifo_store[19][3] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_02924_));
 sky130_fd_sc_hd__mux4_1 _13843_ (.A0(\fifo0.fifo_store[20][3] ),
    .A1(\fifo0.fifo_store[21][3] ),
    .A2(\fifo0.fifo_store[22][3] ),
    .A3(\fifo0.fifo_store[23][3] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _13844_ (.A0(_02924_),
    .A1(_02925_),
    .S(_06565_),
    .X(_02926_));
 sky130_fd_sc_hd__mux4_1 _13845_ (.A0(\fifo0.fifo_store[28][3] ),
    .A1(\fifo0.fifo_store[29][3] ),
    .A2(\fifo0.fifo_store[30][3] ),
    .A3(\fifo0.fifo_store[31][3] ),
    .S0(_06451_),
    .S1(_06453_),
    .X(_02927_));
 sky130_fd_sc_hd__or2_1 _13846_ (.A(_06502_),
    .B(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__mux4_1 _13847_ (.A0(\fifo0.fifo_store[24][3] ),
    .A1(\fifo0.fifo_store[25][3] ),
    .A2(\fifo0.fifo_store[26][3] ),
    .A3(\fifo0.fifo_store[27][3] ),
    .S0(_06600_),
    .S1(_06555_),
    .X(_02929_));
 sky130_fd_sc_hd__o21a_1 _13848_ (.A1(_06599_),
    .A2(_02929_),
    .B1(_06571_),
    .X(_02930_));
 sky130_fd_sc_hd__a221o_1 _13849_ (.A1(_06552_),
    .A2(_02926_),
    .B1(_02928_),
    .B2(_02930_),
    .C1(_06494_),
    .X(_02931_));
 sky130_fd_sc_hd__o311a_1 _13850_ (.A1(_06409_),
    .A2(_02919_),
    .A3(_02923_),
    .B1(_02931_),
    .C1(_06575_),
    .X(_02932_));
 sky130_fd_sc_hd__mux4_1 _13851_ (.A0(\fifo0.fifo_store[36][3] ),
    .A1(\fifo0.fifo_store[37][3] ),
    .A2(\fifo0.fifo_store[38][3] ),
    .A3(\fifo0.fifo_store[39][3] ),
    .S0(_06452_),
    .S1(_06454_),
    .X(_02933_));
 sky130_fd_sc_hd__mux4_1 _13852_ (.A0(\fifo0.fifo_store[32][3] ),
    .A1(\fifo0.fifo_store[33][3] ),
    .A2(\fifo0.fifo_store[34][3] ),
    .A3(\fifo0.fifo_store[35][3] ),
    .S0(_06977_),
    .S1(_06437_),
    .X(_02934_));
 sky130_fd_sc_hd__or2_1 _13853_ (.A(_06441_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__o211a_1 _13854_ (.A1(_07355_),
    .A2(_02933_),
    .B1(_02935_),
    .C1(_06468_),
    .X(_02936_));
 sky130_fd_sc_hd__mux4_1 _13855_ (.A0(\fifo0.fifo_store[40][3] ),
    .A1(\fifo0.fifo_store[41][3] ),
    .A2(\fifo0.fifo_store[42][3] ),
    .A3(\fifo0.fifo_store[43][3] ),
    .S0(_06951_),
    .S1(_06556_),
    .X(_02937_));
 sky130_fd_sc_hd__or2b_1 _13856_ (.A(\fifo0.fifo_store[47][3] ),
    .B_N(_07097_),
    .X(_02938_));
 sky130_fd_sc_hd__o21a_1 _13857_ (.A1(_07097_),
    .A2(\fifo0.fifo_store[46][3] ),
    .B1(_06421_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _13858_ (.A0(\fifo0.fifo_store[44][3] ),
    .A1(\fifo0.fifo_store[45][3] ),
    .S(_06946_),
    .X(_02940_));
 sky130_fd_sc_hd__a221o_1 _13859_ (.A1(_02938_),
    .A2(_02939_),
    .B1(_02940_),
    .B2(_06425_),
    .C1(_06502_),
    .X(_02941_));
 sky130_fd_sc_hd__o211a_1 _13860_ (.A1(_06554_),
    .A2(_02937_),
    .B1(_02941_),
    .C1(_06463_),
    .X(_02942_));
 sky130_fd_sc_hd__mux4_1 _13861_ (.A0(\fifo0.fifo_store[48][3] ),
    .A1(\fifo0.fifo_store[49][3] ),
    .A2(\fifo0.fifo_store[50][3] ),
    .A3(\fifo0.fifo_store[51][3] ),
    .S0(_06591_),
    .S1(_06592_),
    .X(_02943_));
 sky130_fd_sc_hd__mux4_1 _13862_ (.A0(\fifo0.fifo_store[52][3] ),
    .A1(\fifo0.fifo_store[53][3] ),
    .A2(\fifo0.fifo_store[54][3] ),
    .A3(\fifo0.fifo_store[55][3] ),
    .S0(_06977_),
    .S1(_06437_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _13863_ (.A0(_02943_),
    .A1(_02944_),
    .S(_06474_),
    .X(_02945_));
 sky130_fd_sc_hd__mux4_1 _13864_ (.A0(\fifo0.fifo_store[60][3] ),
    .A1(\fifo0.fifo_store[61][3] ),
    .A2(\fifo0.fifo_store[62][3] ),
    .A3(\fifo0.fifo_store[63][3] ),
    .S0(_07017_),
    .S1(_07391_),
    .X(_02946_));
 sky130_fd_sc_hd__or2_1 _13865_ (.A(_07371_),
    .B(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__mux4_1 _13866_ (.A0(\fifo0.fifo_store[56][3] ),
    .A1(\fifo0.fifo_store[57][3] ),
    .A2(\fifo0.fifo_store[58][3] ),
    .A3(\fifo0.fifo_store[59][3] ),
    .S0(_06693_),
    .S1(_06579_),
    .X(_02948_));
 sky130_fd_sc_hd__o21a_1 _13867_ (.A1(_06624_),
    .A2(_02948_),
    .B1(_07219_),
    .X(_02949_));
 sky130_fd_sc_hd__a221o_2 _13868_ (.A1(_06793_),
    .A2(_02945_),
    .B1(_02947_),
    .B2(_02949_),
    .C1(_06494_),
    .X(_02950_));
 sky130_fd_sc_hd__o311a_1 _13869_ (.A1(_06409_),
    .A2(_02936_),
    .A3(_02942_),
    .B1(_06465_),
    .C1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__o31a_1 _13870_ (.A1(_06992_),
    .A2(_02932_),
    .A3(_02951_),
    .B1(_06606_),
    .X(_02952_));
 sky130_fd_sc_hd__a211oi_1 _13871_ (.A1(_06370_),
    .A2(_06757_),
    .B1(_06392_),
    .C1(_06359_),
    .Y(_02953_));
 sky130_fd_sc_hd__inv_2 _13872_ (.A(_06775_),
    .Y(_02954_));
 sky130_fd_sc_hd__a2bb2o_1 _13873_ (.A1_N(_06891_),
    .A2_N(_02954_),
    .B1(_06910_),
    .B2(_06386_),
    .X(_02955_));
 sky130_fd_sc_hd__or2_1 _13874_ (.A(_06747_),
    .B(_02665_),
    .X(_02956_));
 sky130_fd_sc_hd__o21ai_1 _13875_ (.A1(_02953_),
    .A2(_02955_),
    .B1(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__o311a_1 _13876_ (.A1(_06919_),
    .A2(_02953_),
    .A3(_02955_),
    .B1(_02957_),
    .C1(_06918_),
    .X(_02958_));
 sky130_fd_sc_hd__a211o_1 _13877_ (.A1(_02913_),
    .A2(_02952_),
    .B1(_06353_),
    .C1(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__a21o_1 _13878_ (.A1(_02862_),
    .A2(_02959_),
    .B1(net31),
    .X(_02960_));
 sky130_fd_sc_hd__o21a_1 _13879_ (.A1(_07315_),
    .A2(_02764_),
    .B1(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__mux4_1 _13880_ (.A0(_07167_),
    .A1(_02771_),
    .A2(_02772_),
    .A3(_02961_),
    .S0(_07326_),
    .S1(_07314_),
    .X(_02962_));
 sky130_fd_sc_hd__and2_1 _13881_ (.A(_07331_),
    .B(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__nand2_1 _13882_ (.A(\dsmod0.accu1[3] ),
    .B(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__mux4_1 _13883_ (.A0(_02171_),
    .A1(_02370_),
    .A2(_02573_),
    .A3(_02763_),
    .S0(_07164_),
    .S1(_07165_),
    .X(_02965_));
 sky130_fd_sc_hd__or2_1 _13884_ (.A(_07326_),
    .B(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__a21oi_1 _13885_ (.A1(_02913_),
    .A2(_02952_),
    .B1(_02958_),
    .Y(_02967_));
 sky130_fd_sc_hd__or2_1 _13886_ (.A(_02205_),
    .B(\fifo0.fifo_store[103][2] ),
    .X(_02968_));
 sky130_fd_sc_hd__o21a_1 _13887_ (.A1(_02871_),
    .A2(\fifo0.fifo_store[102][2] ),
    .B1(_06438_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _13888_ (.A0(\fifo0.fifo_store[100][2] ),
    .A1(\fifo0.fifo_store[101][2] ),
    .S(_06951_),
    .X(_02970_));
 sky130_fd_sc_hd__a221o_1 _13889_ (.A1(_02968_),
    .A2(_02969_),
    .B1(_02970_),
    .B2(_06954_),
    .C1(_06945_),
    .X(_02971_));
 sky130_fd_sc_hd__mux4_1 _13890_ (.A0(\fifo0.fifo_store[96][2] ),
    .A1(\fifo0.fifo_store[97][2] ),
    .A2(\fifo0.fifo_store[98][2] ),
    .A3(\fifo0.fifo_store[99][2] ),
    .S0(_07067_),
    .S1(_06971_),
    .X(_02972_));
 sky130_fd_sc_hd__or2_1 _13891_ (.A(_07066_),
    .B(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__mux4_2 _13892_ (.A0(\fifo0.fifo_store[104][2] ),
    .A1(\fifo0.fifo_store[105][2] ),
    .A2(\fifo0.fifo_store[106][2] ),
    .A3(\fifo0.fifo_store[107][2] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_02974_));
 sky130_fd_sc_hd__mux4_1 _13893_ (.A0(\fifo0.fifo_store[108][2] ),
    .A1(\fifo0.fifo_store[109][2] ),
    .A2(\fifo0.fifo_store[110][2] ),
    .A3(\fifo0.fifo_store[111][2] ),
    .S0(_07008_),
    .S1(_06725_),
    .X(_02975_));
 sky130_fd_sc_hd__or2_1 _13894_ (.A(_06709_),
    .B(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__o211a_1 _13895_ (.A1(_07066_),
    .A2(_02974_),
    .B1(_02976_),
    .C1(_07094_),
    .X(_02977_));
 sky130_fd_sc_hd__a311o_1 _13896_ (.A1(_06939_),
    .A2(_02971_),
    .A3(_02973_),
    .B1(_02977_),
    .C1(_06409_),
    .X(_02978_));
 sky130_fd_sc_hd__mux4_1 _13897_ (.A0(\fifo0.fifo_store[112][2] ),
    .A1(\fifo0.fifo_store[113][2] ),
    .A2(\fifo0.fifo_store[114][2] ),
    .A3(\fifo0.fifo_store[115][2] ),
    .S0(_06416_),
    .S1(_06691_),
    .X(_02979_));
 sky130_fd_sc_hd__mux4_1 _13898_ (.A0(\fifo0.fifo_store[116][2] ),
    .A1(\fifo0.fifo_store[117][2] ),
    .A2(\fifo0.fifo_store[118][2] ),
    .A3(\fifo0.fifo_store[119][2] ),
    .S0(_07001_),
    .S1(_06691_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _13899_ (.A0(_02979_),
    .A1(_02980_),
    .S(_06824_),
    .X(_02981_));
 sky130_fd_sc_hd__mux4_1 _13900_ (.A0(\fifo0.fifo_store[124][2] ),
    .A1(\fifo0.fifo_store[125][2] ),
    .A2(\fifo0.fifo_store[126][2] ),
    .A3(\fifo0.fifo_store[127][2] ),
    .S0(_06508_),
    .S1(_06996_),
    .X(_02982_));
 sky130_fd_sc_hd__or2_1 _13901_ (.A(_07071_),
    .B(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__mux4_2 _13902_ (.A0(\fifo0.fifo_store[120][2] ),
    .A1(\fifo0.fifo_store[121][2] ),
    .A2(\fifo0.fifo_store[122][2] ),
    .A3(\fifo0.fifo_store[123][2] ),
    .S0(_07097_),
    .S1(_07099_),
    .X(_02984_));
 sky130_fd_sc_hd__o21a_1 _13903_ (.A1(_07096_),
    .A2(_02984_),
    .B1(_07094_),
    .X(_02985_));
 sky130_fd_sc_hd__a221o_1 _13904_ (.A1(_06939_),
    .A2(_02981_),
    .B1(_02983_),
    .B2(_02985_),
    .C1(_07085_),
    .X(_02986_));
 sky130_fd_sc_hd__mux4_2 _13905_ (.A0(\fifo0.fifo_store[84][2] ),
    .A1(\fifo0.fifo_store[85][2] ),
    .A2(\fifo0.fifo_store[86][2] ),
    .A3(\fifo0.fifo_store[87][2] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_02987_));
 sky130_fd_sc_hd__mux4_1 _13906_ (.A0(\fifo0.fifo_store[80][2] ),
    .A1(\fifo0.fifo_store[81][2] ),
    .A2(\fifo0.fifo_store[82][2] ),
    .A3(\fifo0.fifo_store[83][2] ),
    .S0(_07008_),
    .S1(_06725_),
    .X(_02988_));
 sky130_fd_sc_hd__or2_1 _13907_ (.A(_06565_),
    .B(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__o211a_1 _13908_ (.A1(_07071_),
    .A2(_02987_),
    .B1(_02989_),
    .C1(_07107_),
    .X(_02990_));
 sky130_fd_sc_hd__buf_8 _13909_ (.A(_07209_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _13910_ (.A0(\fifo0.fifo_store[94][2] ),
    .A1(\fifo0.fifo_store[95][2] ),
    .S(_07079_),
    .X(_02992_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_02991_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__mux2_1 _13912_ (.A0(\fifo0.fifo_store[92][2] ),
    .A1(\fifo0.fifo_store[93][2] ),
    .S(_06951_),
    .X(_02994_));
 sky130_fd_sc_hd__a21oi_1 _13913_ (.A1(_06954_),
    .A2(_02994_),
    .B1(_07071_),
    .Y(_02995_));
 sky130_fd_sc_hd__mux4_2 _13914_ (.A0(\fifo0.fifo_store[88][2] ),
    .A1(\fifo0.fifo_store[89][2] ),
    .A2(\fifo0.fifo_store[90][2] ),
    .A3(\fifo0.fifo_store[91][2] ),
    .S0(_06576_),
    .S1(_07073_),
    .X(_02996_));
 sky130_fd_sc_hd__o21ai_1 _13915_ (.A1(_07096_),
    .A2(_02996_),
    .B1(_07094_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21oi_1 _13916_ (.A1(_02993_),
    .A2(_02995_),
    .B1(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__mux4_2 _13917_ (.A0(\fifo0.fifo_store[64][2] ),
    .A1(\fifo0.fifo_store[65][2] ),
    .A2(\fifo0.fifo_store[66][2] ),
    .A3(\fifo0.fifo_store[67][2] ),
    .S0(_06710_),
    .S1(_06984_),
    .X(_02999_));
 sky130_fd_sc_hd__mux4_1 _13918_ (.A0(\fifo0.fifo_store[68][2] ),
    .A1(\fifo0.fifo_store[69][2] ),
    .A2(\fifo0.fifo_store[70][2] ),
    .A3(\fifo0.fifo_store[71][2] ),
    .S0(_06415_),
    .S1(_06984_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _13919_ (.A0(_02999_),
    .A1(_03000_),
    .S(_06730_),
    .X(_03001_));
 sky130_fd_sc_hd__mux4_1 _13920_ (.A0(\fifo0.fifo_store[76][2] ),
    .A1(\fifo0.fifo_store[77][2] ),
    .A2(\fifo0.fifo_store[78][2] ),
    .A3(\fifo0.fifo_store[79][2] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_03002_));
 sky130_fd_sc_hd__or2_1 _13921_ (.A(_07070_),
    .B(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__mux4_1 _13922_ (.A0(\fifo0.fifo_store[72][2] ),
    .A1(\fifo0.fifo_store[73][2] ),
    .A2(\fifo0.fifo_store[74][2] ),
    .A3(\fifo0.fifo_store[75][2] ),
    .S0(_06434_),
    .S1(_07098_),
    .X(_03004_));
 sky130_fd_sc_hd__o21a_1 _13923_ (.A1(_06441_),
    .A2(_03004_),
    .B1(_06713_),
    .X(_03005_));
 sky130_fd_sc_hd__a221o_1 _13924_ (.A1(_07107_),
    .A2(_03001_),
    .B1(_03003_),
    .B2(_03005_),
    .C1(_06408_),
    .X(_03006_));
 sky130_fd_sc_hd__o311a_1 _13925_ (.A1(_07085_),
    .A2(_02990_),
    .A3(_02998_),
    .B1(_03006_),
    .C1(_06498_),
    .X(_03007_));
 sky130_fd_sc_hd__a311o_4 _13926_ (.A1(_06792_),
    .A2(_02978_),
    .A3(_02986_),
    .B1(_03007_),
    .C1(_06965_),
    .X(_03008_));
 sky130_fd_sc_hd__or2_1 _13927_ (.A(_06416_),
    .B(\fifo0.fifo_store[38][2] ),
    .X(_03009_));
 sky130_fd_sc_hd__o211a_1 _13928_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[39][2] ),
    .B1(_03009_),
    .C1(_06422_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _13929_ (.A0(\fifo0.fifo_store[36][2] ),
    .A1(\fifo0.fifo_store[37][2] ),
    .S(_07227_),
    .X(_03011_));
 sky130_fd_sc_hd__a21o_1 _13930_ (.A1(_06425_),
    .A2(_03011_),
    .B1(_06517_),
    .X(_03012_));
 sky130_fd_sc_hd__mux4_1 _13931_ (.A0(\fifo0.fifo_store[32][2] ),
    .A1(\fifo0.fifo_store[33][2] ),
    .A2(\fifo0.fifo_store[34][2] ),
    .A3(\fifo0.fifo_store[35][2] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_03013_));
 sky130_fd_sc_hd__o221a_1 _13932_ (.A1(_03010_),
    .A2(_03012_),
    .B1(_03013_),
    .B2(_06442_),
    .C1(_06552_),
    .X(_03014_));
 sky130_fd_sc_hd__mux4_1 _13933_ (.A0(\fifo0.fifo_store[40][2] ),
    .A1(\fifo0.fifo_store[41][2] ),
    .A2(\fifo0.fifo_store[42][2] ),
    .A3(\fifo0.fifo_store[43][2] ),
    .S0(_06951_),
    .S1(_06556_),
    .X(_03015_));
 sky130_fd_sc_hd__mux4_1 _13934_ (.A0(\fifo0.fifo_store[44][2] ),
    .A1(\fifo0.fifo_store[45][2] ),
    .A2(\fifo0.fifo_store[46][2] ),
    .A3(\fifo0.fifo_store[47][2] ),
    .S0(_06795_),
    .S1(_06453_),
    .X(_03016_));
 sky130_fd_sc_hd__or2_1 _13935_ (.A(_06502_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _13936_ (.A1(_06554_),
    .A2(_03015_),
    .B1(_03017_),
    .C1(_06463_),
    .X(_03018_));
 sky130_fd_sc_hd__mux4_1 _13937_ (.A0(\fifo0.fifo_store[48][2] ),
    .A1(\fifo0.fifo_store[49][2] ),
    .A2(\fifo0.fifo_store[50][2] ),
    .A3(\fifo0.fifo_store[51][2] ),
    .S0(_02265_),
    .S1(_06437_),
    .X(_03019_));
 sky130_fd_sc_hd__mux4_1 _13938_ (.A0(\fifo0.fifo_store[52][2] ),
    .A1(\fifo0.fifo_store[53][2] ),
    .A2(\fifo0.fifo_store[54][2] ),
    .A3(\fifo0.fifo_store[55][2] ),
    .S0(_02265_),
    .S1(_06471_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _13939_ (.A0(_03019_),
    .A1(_03020_),
    .S(_06474_),
    .X(_03021_));
 sky130_fd_sc_hd__mux4_2 _13940_ (.A0(\fifo0.fifo_store[60][2] ),
    .A1(\fifo0.fifo_store[61][2] ),
    .A2(\fifo0.fifo_store[62][2] ),
    .A3(\fifo0.fifo_store[63][2] ),
    .S0(_06569_),
    .S1(_06481_),
    .X(_03022_));
 sky130_fd_sc_hd__or2_1 _13941_ (.A(_06477_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__mux4_1 _13942_ (.A0(\fifo0.fifo_store[56][2] ),
    .A1(\fifo0.fifo_store[57][2] ),
    .A2(\fifo0.fifo_store[58][2] ),
    .A3(\fifo0.fifo_store[59][2] ),
    .S0(_06625_),
    .S1(_06489_),
    .X(_03024_));
 sky130_fd_sc_hd__o21a_1 _13943_ (.A1(_06624_),
    .A2(_03024_),
    .B1(_07219_),
    .X(_03025_));
 sky130_fd_sc_hd__a221o_2 _13944_ (.A1(_06468_),
    .A2(_03021_),
    .B1(_03023_),
    .B2(_03025_),
    .C1(_06494_),
    .X(_03026_));
 sky130_fd_sc_hd__o311a_1 _13945_ (.A1(_06409_),
    .A2(_03014_),
    .A3(_03018_),
    .B1(_06465_),
    .C1(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__mux4_1 _13946_ (.A0(\fifo0.fifo_store[0][2] ),
    .A1(\fifo0.fifo_store[1][2] ),
    .A2(\fifo0.fifo_store[2][2] ),
    .A3(\fifo0.fifo_store[3][2] ),
    .S0(_06977_),
    .S1(_06592_),
    .X(_03028_));
 sky130_fd_sc_hd__or2_1 _13947_ (.A(_06448_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__mux4_1 _13948_ (.A0(\fifo0.fifo_store[4][2] ),
    .A1(\fifo0.fifo_store[5][2] ),
    .A2(\fifo0.fifo_store[6][2] ),
    .A3(\fifo0.fifo_store[7][2] ),
    .S0(_06503_),
    .S1(_06504_),
    .X(_03030_));
 sky130_fd_sc_hd__o21a_1 _13949_ (.A1(_06502_),
    .A2(_03030_),
    .B1(_06444_),
    .X(_03031_));
 sky130_fd_sc_hd__or2b_1 _13950_ (.A(\fifo0.fifo_store[15][2] ),
    .B_N(_06508_),
    .X(_03032_));
 sky130_fd_sc_hd__o21a_1 _13951_ (.A1(_06508_),
    .A2(\fifo0.fifo_store[14][2] ),
    .B1(_06511_),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _13952_ (.A0(\fifo0.fifo_store[12][2] ),
    .A1(\fifo0.fifo_store[13][2] ),
    .S(_06959_),
    .X(_03034_));
 sky130_fd_sc_hd__a221o_1 _13953_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03034_),
    .B2(_06516_),
    .C1(_06456_),
    .X(_03035_));
 sky130_fd_sc_hd__mux4_2 _13954_ (.A0(\fifo0.fifo_store[8][2] ),
    .A1(\fifo0.fifo_store[9][2] ),
    .A2(\fifo0.fifo_store[10][2] ),
    .A3(\fifo0.fifo_store[11][2] ),
    .S0(_06600_),
    .S1(_06555_),
    .X(_03036_));
 sky130_fd_sc_hd__o21a_1 _13955_ (.A1(_06599_),
    .A2(_03036_),
    .B1(_06571_),
    .X(_03037_));
 sky130_fd_sc_hd__a221o_1 _13956_ (.A1(_03029_),
    .A2(_03031_),
    .B1(_03035_),
    .B2(_03037_),
    .C1(_06408_),
    .X(_03038_));
 sky130_fd_sc_hd__mux4_1 _13957_ (.A0(\fifo0.fifo_store[16][2] ),
    .A1(\fifo0.fifo_store[17][2] ),
    .A2(\fifo0.fifo_store[18][2] ),
    .A3(\fifo0.fifo_store[19][2] ),
    .S0(_06645_),
    .S1(_07111_),
    .X(_03039_));
 sky130_fd_sc_hd__mux4_1 _13958_ (.A0(\fifo0.fifo_store[20][2] ),
    .A1(\fifo0.fifo_store[21][2] ),
    .A2(\fifo0.fifo_store[22][2] ),
    .A3(\fifo0.fifo_store[23][2] ),
    .S0(_06527_),
    .S1(_06528_),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _13959_ (.A0(_03039_),
    .A1(_03040_),
    .S(_06531_),
    .X(_03041_));
 sky130_fd_sc_hd__mux4_1 _13960_ (.A0(\fifo0.fifo_store[28][2] ),
    .A1(\fifo0.fifo_store[29][2] ),
    .A2(\fifo0.fifo_store[30][2] ),
    .A3(\fifo0.fifo_store[31][2] ),
    .S0(_06457_),
    .S1(_06458_),
    .X(_03042_));
 sky130_fd_sc_hd__or2_1 _13961_ (.A(_06456_),
    .B(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__mux4_2 _13962_ (.A0(\fifo0.fifo_store[24][2] ),
    .A1(\fifo0.fifo_store[25][2] ),
    .A2(\fifo0.fifo_store[26][2] ),
    .A3(\fifo0.fifo_store[27][2] ),
    .S0(_06521_),
    .S1(_06523_),
    .X(_03044_));
 sky130_fd_sc_hd__o21a_1 _13963_ (.A1(_06519_),
    .A2(_03044_),
    .B1(_06571_),
    .X(_03045_));
 sky130_fd_sc_hd__a221o_1 _13964_ (.A1(_06445_),
    .A2(_03041_),
    .B1(_03043_),
    .B2(_03045_),
    .C1(_06539_),
    .X(_03046_));
 sky130_fd_sc_hd__a31o_1 _13965_ (.A1(_06498_),
    .A2(_03038_),
    .A3(_03046_),
    .B1(_00006_),
    .X(_03047_));
 sky130_fd_sc_hd__o21a_1 _13966_ (.A1(_03027_),
    .A2(_03047_),
    .B1(_06606_),
    .X(_03048_));
 sky130_fd_sc_hd__o32a_1 _13967_ (.A1(_06374_),
    .A2(_02954_),
    .A3(_06400_),
    .B1(_07198_),
    .B2(_06891_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _13968_ (.A0(_06769_),
    .A1(_02956_),
    .S(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__o2bb2a_1 _13969_ (.A1_N(_03008_),
    .A2_N(_03048_),
    .B1(_06611_),
    .B2(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _13970_ (.A0(_02967_),
    .A1(_03051_),
    .S(_07164_),
    .X(_03052_));
 sky130_fd_sc_hd__a211o_1 _13971_ (.A1(_06611_),
    .A2(_02852_),
    .B1(_02861_),
    .C1(_06353_),
    .X(_03053_));
 sky130_fd_sc_hd__o21ai_1 _13972_ (.A1(_07322_),
    .A2(_02668_),
    .B1(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__nor2_1 _13973_ (.A(_07165_),
    .B(net32),
    .Y(_03055_));
 sky130_fd_sc_hd__a221oi_4 _13974_ (.A1(_07171_),
    .A2(_03052_),
    .B1(_03054_),
    .B2(_03055_),
    .C1(_06354_),
    .Y(_03056_));
 sky130_fd_sc_hd__a32oi_4 _13975_ (.A1(_06354_),
    .A2(_07320_),
    .A3(_07327_),
    .B1(_02966_),
    .B2(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__nor2_1 _13976_ (.A(_06356_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _13977_ (.A(\dsmod0.accu1[2] ),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__and3b_1 _13978_ (.A_N(_02665_),
    .B(_06918_),
    .C(_06919_),
    .X(_03060_));
 sky130_fd_sc_hd__buf_4 _13979_ (.A(_07132_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_4 _13980_ (.A(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__buf_4 _13981_ (.A(_07204_),
    .X(_03063_));
 sky130_fd_sc_hd__mux4_1 _13982_ (.A0(\fifo0.fifo_store[28][0] ),
    .A1(\fifo0.fifo_store[29][0] ),
    .A2(\fifo0.fifo_store[30][0] ),
    .A3(\fifo0.fifo_store[31][0] ),
    .S0(_03063_),
    .S1(_02897_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_4 _13983_ (.A(_06442_),
    .X(_03065_));
 sky130_fd_sc_hd__buf_6 _13984_ (.A(_07079_),
    .X(_03066_));
 sky130_fd_sc_hd__mux4_1 _13985_ (.A0(\fifo0.fifo_store[24][0] ),
    .A1(\fifo0.fifo_store[25][0] ),
    .A2(\fifo0.fifo_store[26][0] ),
    .A3(\fifo0.fifo_store[27][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03067_));
 sky130_fd_sc_hd__or2_1 _13986_ (.A(_03065_),
    .B(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__buf_4 _13987_ (.A(_07220_),
    .X(_03069_));
 sky130_fd_sc_hd__o211a_1 _13988_ (.A1(_03062_),
    .A2(_03064_),
    .B1(_03068_),
    .C1(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__or2_1 _13989_ (.A(_03063_),
    .B(\fifo0.fifo_store[22][0] ),
    .X(_03071_));
 sky130_fd_sc_hd__o211a_1 _13990_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[23][0] ),
    .B1(_03071_),
    .C1(_02897_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _13991_ (.A0(\fifo0.fifo_store[20][0] ),
    .A1(\fifo0.fifo_store[21][0] ),
    .S(_03063_),
    .X(_03073_));
 sky130_fd_sc_hd__a21o_1 _13992_ (.A1(_07207_),
    .A2(_03073_),
    .B1(_03062_),
    .X(_03074_));
 sky130_fd_sc_hd__mux4_1 _13993_ (.A0(\fifo0.fifo_store[16][0] ),
    .A1(\fifo0.fifo_store[17][0] ),
    .A2(\fifo0.fifo_store[18][0] ),
    .A3(\fifo0.fifo_store[19][0] ),
    .S0(_03063_),
    .S1(_02897_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_4 _13994_ (.A(_06793_),
    .X(_03076_));
 sky130_fd_sc_hd__o221a_1 _13995_ (.A1(_03072_),
    .A2(_03074_),
    .B1(_03075_),
    .B2(_03065_),
    .C1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__mux4_1 _13996_ (.A0(\fifo0.fifo_store[0][0] ),
    .A1(\fifo0.fifo_store[1][0] ),
    .A2(\fifo0.fifo_store[2][0] ),
    .A3(\fifo0.fifo_store[3][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03078_));
 sky130_fd_sc_hd__or2_1 _13997_ (.A(_03065_),
    .B(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__mux4_1 _13998_ (.A0(\fifo0.fifo_store[4][0] ),
    .A1(\fifo0.fifo_store[5][0] ),
    .A2(\fifo0.fifo_store[6][0] ),
    .A3(\fifo0.fifo_store[7][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03080_));
 sky130_fd_sc_hd__or2_1 _13999_ (.A(_03061_),
    .B(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__buf_8 _14000_ (.A(_02871_),
    .X(_03082_));
 sky130_fd_sc_hd__buf_6 _14001_ (.A(_07205_),
    .X(_03083_));
 sky130_fd_sc_hd__mux4_1 _14002_ (.A0(\fifo0.fifo_store[12][0] ),
    .A1(\fifo0.fifo_store[13][0] ),
    .A2(\fifo0.fifo_store[14][0] ),
    .A3(\fifo0.fifo_store[15][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__mux4_1 _14003_ (.A0(\fifo0.fifo_store[8][0] ),
    .A1(\fifo0.fifo_store[9][0] ),
    .A2(\fifo0.fifo_store[10][0] ),
    .A3(\fifo0.fifo_store[11][0] ),
    .S0(_02871_),
    .S1(_07205_),
    .X(_03085_));
 sky130_fd_sc_hd__or2_1 _14004_ (.A(_02894_),
    .B(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__o211a_1 _14005_ (.A1(_03062_),
    .A2(_03084_),
    .B1(_03086_),
    .C1(_03069_),
    .X(_03087_));
 sky130_fd_sc_hd__a311o_1 _14006_ (.A1(_03076_),
    .A2(_03079_),
    .A3(_03081_),
    .B1(_07202_),
    .C1(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__o311a_1 _14007_ (.A1(_07354_),
    .A2(_03070_),
    .A3(_03077_),
    .B1(_03088_),
    .C1(_06575_),
    .X(_03089_));
 sky130_fd_sc_hd__mux4_1 _14008_ (.A0(\fifo0.fifo_store[56][0] ),
    .A1(\fifo0.fifo_store[57][0] ),
    .A2(\fifo0.fifo_store[58][0] ),
    .A3(\fifo0.fifo_store[59][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03090_));
 sky130_fd_sc_hd__or2_1 _14009_ (.A(_03065_),
    .B(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__or2_1 _14010_ (.A(_02234_),
    .B(\fifo0.fifo_store[63][0] ),
    .X(_03092_));
 sky130_fd_sc_hd__o21a_1 _14011_ (.A1(_03063_),
    .A2(\fifo0.fifo_store[62][0] ),
    .B1(_02897_),
    .X(_03093_));
 sky130_fd_sc_hd__mux2_1 _14012_ (.A0(\fifo0.fifo_store[60][0] ),
    .A1(\fifo0.fifo_store[61][0] ),
    .S(_03082_),
    .X(_03094_));
 sky130_fd_sc_hd__a221o_1 _14013_ (.A1(_03092_),
    .A2(_03093_),
    .B1(_03094_),
    .B2(_07207_),
    .C1(_03061_),
    .X(_03095_));
 sky130_fd_sc_hd__mux4_1 _14014_ (.A0(\fifo0.fifo_store[52][0] ),
    .A1(\fifo0.fifo_store[53][0] ),
    .A2(\fifo0.fifo_store[54][0] ),
    .A3(\fifo0.fifo_store[55][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03096_));
 sky130_fd_sc_hd__mux4_1 _14015_ (.A0(\fifo0.fifo_store[48][0] ),
    .A1(\fifo0.fifo_store[49][0] ),
    .A2(\fifo0.fifo_store[50][0] ),
    .A3(\fifo0.fifo_store[51][0] ),
    .S0(_07079_),
    .S1(_07205_),
    .X(_03097_));
 sky130_fd_sc_hd__or2_1 _14016_ (.A(_02894_),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__o211a_1 _14017_ (.A1(_03062_),
    .A2(_03096_),
    .B1(_03098_),
    .C1(_03076_),
    .X(_03099_));
 sky130_fd_sc_hd__a311o_1 _14018_ (.A1(_03069_),
    .A2(_03091_),
    .A3(_03095_),
    .B1(_07354_),
    .C1(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__mux4_1 _14019_ (.A0(\fifo0.fifo_store[32][0] ),
    .A1(\fifo0.fifo_store[33][0] ),
    .A2(\fifo0.fifo_store[34][0] ),
    .A3(\fifo0.fifo_store[35][0] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03101_));
 sky130_fd_sc_hd__mux4_1 _14020_ (.A0(\fifo0.fifo_store[36][0] ),
    .A1(\fifo0.fifo_store[37][0] ),
    .A2(\fifo0.fifo_store[38][0] ),
    .A3(\fifo0.fifo_store[39][0] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _14021_ (.A0(_03101_),
    .A1(_03102_),
    .S(_07203_),
    .X(_03103_));
 sky130_fd_sc_hd__mux4_1 _14022_ (.A0(\fifo0.fifo_store[44][0] ),
    .A1(\fifo0.fifo_store[45][0] ),
    .A2(\fifo0.fifo_store[46][0] ),
    .A3(\fifo0.fifo_store[47][0] ),
    .S0(_03066_),
    .S1(_03083_),
    .X(_03104_));
 sky130_fd_sc_hd__or2_1 _14023_ (.A(_03062_),
    .B(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__mux4_1 _14024_ (.A0(\fifo0.fifo_store[40][0] ),
    .A1(\fifo0.fifo_store[41][0] ),
    .A2(\fifo0.fifo_store[42][0] ),
    .A3(\fifo0.fifo_store[43][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03106_));
 sky130_fd_sc_hd__o21a_1 _14025_ (.A1(_03065_),
    .A2(_03106_),
    .B1(_03069_),
    .X(_03107_));
 sky130_fd_sc_hd__a221o_1 _14026_ (.A1(_03076_),
    .A2(_03103_),
    .B1(_03105_),
    .B2(_03107_),
    .C1(_07202_),
    .X(_03108_));
 sky130_fd_sc_hd__a31o_1 _14027_ (.A1(_06792_),
    .A2(_03100_),
    .A3(_03108_),
    .B1(_06992_),
    .X(_03109_));
 sky130_fd_sc_hd__or2_1 _14028_ (.A(_03063_),
    .B(\fifo0.fifo_store[86][0] ),
    .X(_03110_));
 sky130_fd_sc_hd__o211a_1 _14029_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[87][0] ),
    .B1(_03110_),
    .C1(_02897_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _14030_ (.A0(\fifo0.fifo_store[84][0] ),
    .A1(\fifo0.fifo_store[85][0] ),
    .S(_03063_),
    .X(_03112_));
 sky130_fd_sc_hd__a21o_1 _14031_ (.A1(_07207_),
    .A2(_03112_),
    .B1(_03062_),
    .X(_03113_));
 sky130_fd_sc_hd__mux4_1 _14032_ (.A0(\fifo0.fifo_store[80][0] ),
    .A1(\fifo0.fifo_store[81][0] ),
    .A2(\fifo0.fifo_store[82][0] ),
    .A3(\fifo0.fifo_store[83][0] ),
    .S0(_03063_),
    .S1(_02897_),
    .X(_03114_));
 sky130_fd_sc_hd__o221a_1 _14033_ (.A1(_03111_),
    .A2(_03113_),
    .B1(_03114_),
    .B2(_03065_),
    .C1(_03076_),
    .X(_03115_));
 sky130_fd_sc_hd__mux4_1 _14034_ (.A0(\fifo0.fifo_store[88][0] ),
    .A1(\fifo0.fifo_store[89][0] ),
    .A2(\fifo0.fifo_store[90][0] ),
    .A3(\fifo0.fifo_store[91][0] ),
    .S0(_03063_),
    .S1(_02897_),
    .X(_03116_));
 sky130_fd_sc_hd__mux4_1 _14035_ (.A0(\fifo0.fifo_store[92][0] ),
    .A1(\fifo0.fifo_store[93][0] ),
    .A2(\fifo0.fifo_store[94][0] ),
    .A3(\fifo0.fifo_store[95][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03117_));
 sky130_fd_sc_hd__or2_1 _14036_ (.A(_03062_),
    .B(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__o211a_1 _14037_ (.A1(_03065_),
    .A2(_03116_),
    .B1(_03118_),
    .C1(_03069_),
    .X(_03119_));
 sky130_fd_sc_hd__mux4_1 _14038_ (.A0(\fifo0.fifo_store[64][0] ),
    .A1(\fifo0.fifo_store[65][0] ),
    .A2(\fifo0.fifo_store[66][0] ),
    .A3(\fifo0.fifo_store[67][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03120_));
 sky130_fd_sc_hd__mux4_1 _14039_ (.A0(\fifo0.fifo_store[68][0] ),
    .A1(\fifo0.fifo_store[69][0] ),
    .A2(\fifo0.fifo_store[70][0] ),
    .A3(\fifo0.fifo_store[71][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_1 _14040_ (.A0(_03120_),
    .A1(_03121_),
    .S(_07203_),
    .X(_03122_));
 sky130_fd_sc_hd__mux4_1 _14041_ (.A0(\fifo0.fifo_store[76][0] ),
    .A1(\fifo0.fifo_store[77][0] ),
    .A2(\fifo0.fifo_store[78][0] ),
    .A3(\fifo0.fifo_store[79][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03123_));
 sky130_fd_sc_hd__or2_1 _14042_ (.A(_03062_),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__mux4_1 _14043_ (.A0(\fifo0.fifo_store[72][0] ),
    .A1(\fifo0.fifo_store[73][0] ),
    .A2(\fifo0.fifo_store[74][0] ),
    .A3(\fifo0.fifo_store[75][0] ),
    .S0(_03082_),
    .S1(_02897_),
    .X(_03125_));
 sky130_fd_sc_hd__o21a_1 _14044_ (.A1(_03065_),
    .A2(_03125_),
    .B1(_03069_),
    .X(_03126_));
 sky130_fd_sc_hd__a221o_1 _14045_ (.A1(_03076_),
    .A2(_03122_),
    .B1(_03124_),
    .B2(_03126_),
    .C1(_07202_),
    .X(_03127_));
 sky130_fd_sc_hd__o311a_1 _14046_ (.A1(_07354_),
    .A2(_03115_),
    .A3(_03119_),
    .B1(_03127_),
    .C1(_06575_),
    .X(_03128_));
 sky130_fd_sc_hd__mux4_1 _14047_ (.A0(\fifo0.fifo_store[96][0] ),
    .A1(\fifo0.fifo_store[97][0] ),
    .A2(\fifo0.fifo_store[98][0] ),
    .A3(\fifo0.fifo_store[99][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03129_));
 sky130_fd_sc_hd__or2_1 _14048_ (.A(_03065_),
    .B(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__mux4_1 _14049_ (.A0(\fifo0.fifo_store[100][0] ),
    .A1(\fifo0.fifo_store[101][0] ),
    .A2(\fifo0.fifo_store[102][0] ),
    .A3(\fifo0.fifo_store[103][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03131_));
 sky130_fd_sc_hd__or2_1 _14050_ (.A(_03061_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__mux4_1 _14051_ (.A0(\fifo0.fifo_store[108][0] ),
    .A1(\fifo0.fifo_store[109][0] ),
    .A2(\fifo0.fifo_store[110][0] ),
    .A3(\fifo0.fifo_store[111][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03133_));
 sky130_fd_sc_hd__mux4_1 _14052_ (.A0(\fifo0.fifo_store[104][0] ),
    .A1(\fifo0.fifo_store[105][0] ),
    .A2(\fifo0.fifo_store[106][0] ),
    .A3(\fifo0.fifo_store[107][0] ),
    .S0(_02871_),
    .S1(_07205_),
    .X(_03134_));
 sky130_fd_sc_hd__or2_1 _14053_ (.A(_02894_),
    .B(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__o211a_1 _14054_ (.A1(_03062_),
    .A2(_03133_),
    .B1(_03135_),
    .C1(_03069_),
    .X(_03136_));
 sky130_fd_sc_hd__a311o_1 _14055_ (.A1(_03076_),
    .A2(_03130_),
    .A3(_03132_),
    .B1(_07202_),
    .C1(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__or2_1 _14056_ (.A(_02234_),
    .B(\fifo0.fifo_store[119][0] ),
    .X(_03138_));
 sky130_fd_sc_hd__o21a_1 _14057_ (.A1(_03063_),
    .A2(\fifo0.fifo_store[118][0] ),
    .B1(_02897_),
    .X(_03139_));
 sky130_fd_sc_hd__mux2_1 _14058_ (.A0(\fifo0.fifo_store[116][0] ),
    .A1(\fifo0.fifo_store[117][0] ),
    .S(_03082_),
    .X(_03140_));
 sky130_fd_sc_hd__a221o_1 _14059_ (.A1(_03138_),
    .A2(_03139_),
    .B1(_03140_),
    .B2(_07207_),
    .C1(_03061_),
    .X(_03141_));
 sky130_fd_sc_hd__mux4_1 _14060_ (.A0(\fifo0.fifo_store[112][0] ),
    .A1(\fifo0.fifo_store[113][0] ),
    .A2(\fifo0.fifo_store[114][0] ),
    .A3(\fifo0.fifo_store[115][0] ),
    .S0(_03066_),
    .S1(_02991_),
    .X(_03142_));
 sky130_fd_sc_hd__or2_1 _14061_ (.A(_03065_),
    .B(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__mux4_1 _14062_ (.A0(\fifo0.fifo_store[124][0] ),
    .A1(\fifo0.fifo_store[125][0] ),
    .A2(\fifo0.fifo_store[126][0] ),
    .A3(\fifo0.fifo_store[127][0] ),
    .S0(_03082_),
    .S1(_03083_),
    .X(_03144_));
 sky130_fd_sc_hd__mux4_2 _14063_ (.A0(\fifo0.fifo_store[120][0] ),
    .A1(\fifo0.fifo_store[121][0] ),
    .A2(\fifo0.fifo_store[122][0] ),
    .A3(\fifo0.fifo_store[123][0] ),
    .S0(_02871_),
    .S1(_07205_),
    .X(_03145_));
 sky130_fd_sc_hd__or2_1 _14064_ (.A(_02894_),
    .B(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__o211a_1 _14065_ (.A1(_03062_),
    .A2(_03144_),
    .B1(_03146_),
    .C1(_03069_),
    .X(_03147_));
 sky130_fd_sc_hd__a311o_1 _14066_ (.A1(_03076_),
    .A2(_03141_),
    .A3(_03143_),
    .B1(_07354_),
    .C1(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__a31o_1 _14067_ (.A1(_06792_),
    .A2(_03137_),
    .A3(_03148_),
    .B1(_06965_),
    .X(_03149_));
 sky130_fd_sc_hd__o221a_1 _14068_ (.A1(_03089_),
    .A2(_03109_),
    .B1(_03128_),
    .B2(_03149_),
    .C1(_06611_),
    .X(_03150_));
 sky130_fd_sc_hd__o21ai_1 _14069_ (.A1(_03060_),
    .A2(_03150_),
    .B1(_07322_),
    .Y(_03151_));
 sky130_fd_sc_hd__mux4_1 _14070_ (.A0(\fifo0.fifo_store[28][1] ),
    .A1(\fifo0.fifo_store[29][1] ),
    .A2(\fifo0.fifo_store[30][1] ),
    .A3(\fifo0.fifo_store[31][1] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03152_));
 sky130_fd_sc_hd__mux4_1 _14071_ (.A0(\fifo0.fifo_store[24][1] ),
    .A1(\fifo0.fifo_store[25][1] ),
    .A2(\fifo0.fifo_store[26][1] ),
    .A3(\fifo0.fifo_store[27][1] ),
    .S0(_06951_),
    .S1(_02879_),
    .X(_03153_));
 sky130_fd_sc_hd__or2_1 _14072_ (.A(_06554_),
    .B(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o211a_1 _14073_ (.A1(_03061_),
    .A2(_03152_),
    .B1(_03154_),
    .C1(_03069_),
    .X(_03155_));
 sky130_fd_sc_hd__or2_1 _14074_ (.A(_07204_),
    .B(\fifo0.fifo_store[22][1] ),
    .X(_03156_));
 sky130_fd_sc_hd__o211a_1 _14075_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[23][1] ),
    .B1(_03156_),
    .C1(_03083_),
    .X(_03157_));
 sky130_fd_sc_hd__mux2_1 _14076_ (.A0(\fifo0.fifo_store[20][1] ),
    .A1(\fifo0.fifo_store[21][1] ),
    .S(_07204_),
    .X(_03158_));
 sky130_fd_sc_hd__a21o_1 _14077_ (.A1(_07207_),
    .A2(_03158_),
    .B1(_02866_),
    .X(_03159_));
 sky130_fd_sc_hd__mux4_1 _14078_ (.A0(\fifo0.fifo_store[16][1] ),
    .A1(\fifo0.fifo_store[17][1] ),
    .A2(\fifo0.fifo_store[18][1] ),
    .A3(\fifo0.fifo_store[19][1] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03160_));
 sky130_fd_sc_hd__o221a_1 _14079_ (.A1(_03157_),
    .A2(_03159_),
    .B1(_03160_),
    .B2(_07203_),
    .C1(_03076_),
    .X(_03161_));
 sky130_fd_sc_hd__mux4_2 _14080_ (.A0(\fifo0.fifo_store[8][1] ),
    .A1(\fifo0.fifo_store[9][1] ),
    .A2(\fifo0.fifo_store[10][1] ),
    .A3(\fifo0.fifo_store[11][1] ),
    .S0(_02878_),
    .S1(_07257_),
    .X(_03162_));
 sky130_fd_sc_hd__or2_1 _14081_ (.A(_06554_),
    .B(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__mux4_1 _14082_ (.A0(\fifo0.fifo_store[12][1] ),
    .A1(\fifo0.fifo_store[13][1] ),
    .A2(\fifo0.fifo_store[14][1] ),
    .A3(\fifo0.fifo_store[15][1] ),
    .S0(_07079_),
    .S1(_07209_),
    .X(_03164_));
 sky130_fd_sc_hd__o21a_1 _14083_ (.A1(_03061_),
    .A2(_03164_),
    .B1(_07220_),
    .X(_03165_));
 sky130_fd_sc_hd__mux4_1 _14084_ (.A0(\fifo0.fifo_store[4][1] ),
    .A1(\fifo0.fifo_store[5][1] ),
    .A2(\fifo0.fifo_store[6][1] ),
    .A3(\fifo0.fifo_store[7][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03166_));
 sky130_fd_sc_hd__or2_1 _14085_ (.A(_02866_),
    .B(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__mux4_1 _14086_ (.A0(\fifo0.fifo_store[0][1] ),
    .A1(\fifo0.fifo_store[1][1] ),
    .A2(\fifo0.fifo_store[2][1] ),
    .A3(\fifo0.fifo_store[3][1] ),
    .S0(_07079_),
    .S1(_07209_),
    .X(_03168_));
 sky130_fd_sc_hd__o21a_1 _14087_ (.A1(_02894_),
    .A2(_03168_),
    .B1(_06793_),
    .X(_03169_));
 sky130_fd_sc_hd__a221o_1 _14088_ (.A1(_03163_),
    .A2(_03165_),
    .B1(_03167_),
    .B2(_03169_),
    .C1(_07202_),
    .X(_03170_));
 sky130_fd_sc_hd__o311a_1 _14089_ (.A1(_07354_),
    .A2(_03155_),
    .A3(_03161_),
    .B1(_03170_),
    .C1(_06575_),
    .X(_03171_));
 sky130_fd_sc_hd__mux4_1 _14090_ (.A0(\fifo0.fifo_store[48][1] ),
    .A1(\fifo0.fifo_store[49][1] ),
    .A2(\fifo0.fifo_store[50][1] ),
    .A3(\fifo0.fifo_store[51][1] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_03172_));
 sky130_fd_sc_hd__or2_1 _14091_ (.A(_06554_),
    .B(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__mux4_1 _14092_ (.A0(\fifo0.fifo_store[52][1] ),
    .A1(\fifo0.fifo_store[53][1] ),
    .A2(\fifo0.fifo_store[54][1] ),
    .A3(\fifo0.fifo_store[55][1] ),
    .S0(_02878_),
    .S1(_07257_),
    .X(_03174_));
 sky130_fd_sc_hd__o21a_1 _14093_ (.A1(_02866_),
    .A2(_03174_),
    .B1(_06793_),
    .X(_03175_));
 sky130_fd_sc_hd__or2b_1 _14094_ (.A(\fifo0.fifo_store[63][1] ),
    .B_N(_07204_),
    .X(_03176_));
 sky130_fd_sc_hd__o21a_1 _14095_ (.A1(_07204_),
    .A2(\fifo0.fifo_store[62][1] ),
    .B1(_07209_),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _14096_ (.A0(\fifo0.fifo_store[60][1] ),
    .A1(\fifo0.fifo_store[61][1] ),
    .S(_02871_),
    .X(_03178_));
 sky130_fd_sc_hd__a221o_1 _14097_ (.A1(_03176_),
    .A2(_03177_),
    .B1(_03178_),
    .B2(_07207_),
    .C1(_07355_),
    .X(_03179_));
 sky130_fd_sc_hd__mux4_1 _14098_ (.A0(\fifo0.fifo_store[56][1] ),
    .A1(\fifo0.fifo_store[57][1] ),
    .A2(\fifo0.fifo_store[58][1] ),
    .A3(\fifo0.fifo_store[59][1] ),
    .S0(_02867_),
    .S1(_07257_),
    .X(_03180_));
 sky130_fd_sc_hd__o21a_1 _14099_ (.A1(_02894_),
    .A2(_03180_),
    .B1(_07220_),
    .X(_03181_));
 sky130_fd_sc_hd__a221o_1 _14100_ (.A1(_03173_),
    .A2(_03175_),
    .B1(_03179_),
    .B2(_03181_),
    .C1(_07354_),
    .X(_03182_));
 sky130_fd_sc_hd__mux4_1 _14101_ (.A0(\fifo0.fifo_store[32][1] ),
    .A1(\fifo0.fifo_store[33][1] ),
    .A2(\fifo0.fifo_store[34][1] ),
    .A3(\fifo0.fifo_store[35][1] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_03183_));
 sky130_fd_sc_hd__mux4_1 _14102_ (.A0(\fifo0.fifo_store[36][1] ),
    .A1(\fifo0.fifo_store[37][1] ),
    .A2(\fifo0.fifo_store[38][1] ),
    .A3(\fifo0.fifo_store[39][1] ),
    .S0(_06542_),
    .S1(_06438_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _14103_ (.A0(_03183_),
    .A1(_03184_),
    .S(_07096_),
    .X(_03185_));
 sky130_fd_sc_hd__mux4_1 _14104_ (.A0(\fifo0.fifo_store[44][1] ),
    .A1(\fifo0.fifo_store[45][1] ),
    .A2(\fifo0.fifo_store[46][1] ),
    .A3(\fifo0.fifo_store[47][1] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_03186_));
 sky130_fd_sc_hd__or2_1 _14105_ (.A(_07355_),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__mux4_1 _14106_ (.A0(\fifo0.fifo_store[40][1] ),
    .A1(\fifo0.fifo_store[41][1] ),
    .A2(\fifo0.fifo_store[42][1] ),
    .A3(\fifo0.fifo_store[43][1] ),
    .S0(_02878_),
    .S1(_07257_),
    .X(_03188_));
 sky130_fd_sc_hd__o21a_1 _14107_ (.A1(_06554_),
    .A2(_03188_),
    .B1(_06463_),
    .X(_03189_));
 sky130_fd_sc_hd__a221o_1 _14108_ (.A1(_06939_),
    .A2(_03185_),
    .B1(_03187_),
    .B2(_03189_),
    .C1(_07202_),
    .X(_03190_));
 sky130_fd_sc_hd__a31o_1 _14109_ (.A1(_06792_),
    .A2(_03182_),
    .A3(_03190_),
    .B1(_06992_),
    .X(_03191_));
 sky130_fd_sc_hd__or2_1 _14110_ (.A(_07204_),
    .B(\fifo0.fifo_store[86][1] ),
    .X(_03192_));
 sky130_fd_sc_hd__o211a_1 _14111_ (.A1(_02234_),
    .A2(\fifo0.fifo_store[87][1] ),
    .B1(_03192_),
    .C1(_03083_),
    .X(_03193_));
 sky130_fd_sc_hd__mux2_1 _14112_ (.A0(\fifo0.fifo_store[84][1] ),
    .A1(\fifo0.fifo_store[85][1] ),
    .S(_02871_),
    .X(_03194_));
 sky130_fd_sc_hd__a21o_1 _14113_ (.A1(_07207_),
    .A2(_03194_),
    .B1(_02866_),
    .X(_03195_));
 sky130_fd_sc_hd__mux4_1 _14114_ (.A0(\fifo0.fifo_store[80][1] ),
    .A1(\fifo0.fifo_store[81][1] ),
    .A2(\fifo0.fifo_store[82][1] ),
    .A3(\fifo0.fifo_store[83][1] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03196_));
 sky130_fd_sc_hd__o221a_1 _14115_ (.A1(_03193_),
    .A2(_03195_),
    .B1(_03196_),
    .B2(_07203_),
    .C1(_06939_),
    .X(_03197_));
 sky130_fd_sc_hd__mux4_2 _14116_ (.A0(\fifo0.fifo_store[88][1] ),
    .A1(\fifo0.fifo_store[89][1] ),
    .A2(\fifo0.fifo_store[90][1] ),
    .A3(\fifo0.fifo_store[91][1] ),
    .S0(_02863_),
    .S1(_02864_),
    .X(_03198_));
 sky130_fd_sc_hd__mux4_1 _14117_ (.A0(\fifo0.fifo_store[92][1] ),
    .A1(\fifo0.fifo_store[93][1] ),
    .A2(\fifo0.fifo_store[94][1] ),
    .A3(\fifo0.fifo_store[95][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03199_));
 sky130_fd_sc_hd__or2_1 _14118_ (.A(_02866_),
    .B(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__o211a_1 _14119_ (.A1(_07203_),
    .A2(_03198_),
    .B1(_03200_),
    .C1(_03069_),
    .X(_03201_));
 sky130_fd_sc_hd__mux4_2 _14120_ (.A0(\fifo0.fifo_store[64][1] ),
    .A1(\fifo0.fifo_store[65][1] ),
    .A2(\fifo0.fifo_store[66][1] ),
    .A3(\fifo0.fifo_store[67][1] ),
    .S0(_06951_),
    .S1(_02879_),
    .X(_03202_));
 sky130_fd_sc_hd__mux4_1 _14121_ (.A0(\fifo0.fifo_store[68][1] ),
    .A1(\fifo0.fifo_store[69][1] ),
    .A2(\fifo0.fifo_store[70][1] ),
    .A3(\fifo0.fifo_store[71][1] ),
    .S0(_06951_),
    .S1(_02879_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _14122_ (.A0(_03202_),
    .A1(_03203_),
    .S(_06442_),
    .X(_03204_));
 sky130_fd_sc_hd__mux4_1 _14123_ (.A0(\fifo0.fifo_store[76][1] ),
    .A1(\fifo0.fifo_store[77][1] ),
    .A2(\fifo0.fifo_store[78][1] ),
    .A3(\fifo0.fifo_store[79][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03205_));
 sky130_fd_sc_hd__or2_1 _14124_ (.A(_03061_),
    .B(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__mux4_1 _14125_ (.A0(\fifo0.fifo_store[72][1] ),
    .A1(\fifo0.fifo_store[73][1] ),
    .A2(\fifo0.fifo_store[74][1] ),
    .A3(\fifo0.fifo_store[75][1] ),
    .S0(_07079_),
    .S1(_07209_),
    .X(_03207_));
 sky130_fd_sc_hd__o21a_1 _14126_ (.A1(_02894_),
    .A2(_03207_),
    .B1(_07220_),
    .X(_03208_));
 sky130_fd_sc_hd__a221o_1 _14127_ (.A1(_03076_),
    .A2(_03204_),
    .B1(_03206_),
    .B2(_03208_),
    .C1(_07202_),
    .X(_03209_));
 sky130_fd_sc_hd__o311a_1 _14128_ (.A1(_07354_),
    .A2(_03197_),
    .A3(_03201_),
    .B1(_03209_),
    .C1(_06575_),
    .X(_03210_));
 sky130_fd_sc_hd__mux4_1 _14129_ (.A0(\fifo0.fifo_store[104][1] ),
    .A1(\fifo0.fifo_store[105][1] ),
    .A2(\fifo0.fifo_store[106][1] ),
    .A3(\fifo0.fifo_store[107][1] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_03211_));
 sky130_fd_sc_hd__or2_1 _14130_ (.A(_06554_),
    .B(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__mux4_1 _14131_ (.A0(\fifo0.fifo_store[108][1] ),
    .A1(\fifo0.fifo_store[109][1] ),
    .A2(\fifo0.fifo_store[110][1] ),
    .A3(\fifo0.fifo_store[111][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03213_));
 sky130_fd_sc_hd__o21a_1 _14132_ (.A1(_03061_),
    .A2(_03213_),
    .B1(_07220_),
    .X(_03214_));
 sky130_fd_sc_hd__mux4_1 _14133_ (.A0(\fifo0.fifo_store[100][1] ),
    .A1(\fifo0.fifo_store[101][1] ),
    .A2(\fifo0.fifo_store[102][1] ),
    .A3(\fifo0.fifo_store[103][1] ),
    .S0(_02878_),
    .S1(_07257_),
    .X(_03215_));
 sky130_fd_sc_hd__or2_1 _14134_ (.A(_02866_),
    .B(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__mux4_2 _14135_ (.A0(\fifo0.fifo_store[96][1] ),
    .A1(\fifo0.fifo_store[97][1] ),
    .A2(\fifo0.fifo_store[98][1] ),
    .A3(\fifo0.fifo_store[99][1] ),
    .S0(_02867_),
    .S1(_07209_),
    .X(_03217_));
 sky130_fd_sc_hd__o21a_1 _14136_ (.A1(_02894_),
    .A2(_03217_),
    .B1(_06793_),
    .X(_03218_));
 sky130_fd_sc_hd__a221o_1 _14137_ (.A1(_03212_),
    .A2(_03214_),
    .B1(_03216_),
    .B2(_03218_),
    .C1(_07202_),
    .X(_03219_));
 sky130_fd_sc_hd__mux4_2 _14138_ (.A0(\fifo0.fifo_store[120][1] ),
    .A1(\fifo0.fifo_store[121][1] ),
    .A2(\fifo0.fifo_store[122][1] ),
    .A3(\fifo0.fifo_store[123][1] ),
    .S0(_02878_),
    .S1(_02879_),
    .X(_03220_));
 sky130_fd_sc_hd__or2_1 _14139_ (.A(_06554_),
    .B(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__mux4_1 _14140_ (.A0(\fifo0.fifo_store[124][1] ),
    .A1(\fifo0.fifo_store[125][1] ),
    .A2(\fifo0.fifo_store[126][1] ),
    .A3(\fifo0.fifo_store[127][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03222_));
 sky130_fd_sc_hd__o21a_1 _14141_ (.A1(_03061_),
    .A2(_03222_),
    .B1(_07220_),
    .X(_03223_));
 sky130_fd_sc_hd__or2b_1 _14142_ (.A(\fifo0.fifo_store[119][1] ),
    .B_N(_02863_),
    .X(_03224_));
 sky130_fd_sc_hd__o21a_1 _14143_ (.A1(_02863_),
    .A2(\fifo0.fifo_store[118][1] ),
    .B1(_07205_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _14144_ (.A0(\fifo0.fifo_store[116][1] ),
    .A1(\fifo0.fifo_store[117][1] ),
    .S(_07204_),
    .X(_03226_));
 sky130_fd_sc_hd__a221o_1 _14145_ (.A1(_03224_),
    .A2(_03225_),
    .B1(_03226_),
    .B2(_07207_),
    .C1(_02866_),
    .X(_03227_));
 sky130_fd_sc_hd__mux4_2 _14146_ (.A0(\fifo0.fifo_store[112][1] ),
    .A1(\fifo0.fifo_store[113][1] ),
    .A2(\fifo0.fifo_store[114][1] ),
    .A3(\fifo0.fifo_store[115][1] ),
    .S0(_02867_),
    .S1(_06422_),
    .X(_03228_));
 sky130_fd_sc_hd__o21a_1 _14147_ (.A1(_02894_),
    .A2(_03228_),
    .B1(_06793_),
    .X(_03229_));
 sky130_fd_sc_hd__a221o_1 _14148_ (.A1(_03221_),
    .A2(_03223_),
    .B1(_03227_),
    .B2(_03229_),
    .C1(_07354_),
    .X(_03230_));
 sky130_fd_sc_hd__a31o_1 _14149_ (.A1(_06792_),
    .A2(_03219_),
    .A3(_03230_),
    .B1(_06965_),
    .X(_03231_));
 sky130_fd_sc_hd__o221a_2 _14150_ (.A1(_03171_),
    .A2(_03191_),
    .B1(_03210_),
    .B2(_03231_),
    .C1(_06611_),
    .X(_03232_));
 sky130_fd_sc_hd__nor2_1 _14151_ (.A(_03060_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__o21a_1 _14152_ (.A1(_07322_),
    .A2(_03233_),
    .B1(_07171_),
    .X(_03234_));
 sky130_fd_sc_hd__a22o_1 _14153_ (.A1(_03055_),
    .A2(_03052_),
    .B1(_03151_),
    .B2(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__a21o_1 _14154_ (.A1(_06611_),
    .A2(_02852_),
    .B1(_02861_),
    .X(_03236_));
 sky130_fd_sc_hd__mux4_1 _14155_ (.A0(_02668_),
    .A1(_02573_),
    .A2(_03236_),
    .A3(_02763_),
    .S0(net31),
    .S1(_07322_),
    .X(_03237_));
 sky130_fd_sc_hd__o21ai_1 _14156_ (.A1(_07326_),
    .A2(_03237_),
    .B1(_07314_),
    .Y(_03238_));
 sky130_fd_sc_hd__a2bb2o_1 _14157_ (.A1_N(_03235_),
    .A2_N(_03238_),
    .B1(_06354_),
    .B2(_02376_),
    .X(_03239_));
 sky130_fd_sc_hd__and2_1 _14158_ (.A(_02383_),
    .B(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_1 _14159_ (.A0(_02370_),
    .A1(_02763_),
    .A2(_02573_),
    .A3(_02668_),
    .S0(_07165_),
    .S1(_07322_),
    .X(_03241_));
 sky130_fd_sc_hd__o21ai_1 _14160_ (.A1(_03060_),
    .A2(_03232_),
    .B1(_07322_),
    .Y(_03242_));
 sky130_fd_sc_hd__o211ai_1 _14161_ (.A1(_07322_),
    .A2(_03051_),
    .B1(_03242_),
    .C1(_07171_),
    .Y(_03243_));
 sky130_fd_sc_hd__a21bo_1 _14162_ (.A1(_02862_),
    .A2(_02959_),
    .B1_N(_03055_),
    .X(_03244_));
 sky130_fd_sc_hd__o2111a_1 _14163_ (.A1(_07326_),
    .A2(_03241_),
    .B1(_03243_),
    .C1(_03244_),
    .D1(_07170_),
    .X(_03245_));
 sky130_fd_sc_hd__a211o_1 _14164_ (.A1(_06354_),
    .A2(_02180_),
    .B1(_03245_),
    .C1(_07173_),
    .X(_03246_));
 sky130_fd_sc_hd__a21oi_1 _14165_ (.A1(_07173_),
    .A2(_03233_),
    .B1(_06356_),
    .Y(_03247_));
 sky130_fd_sc_hd__a21o_1 _14166_ (.A1(_03246_),
    .A2(_03247_),
    .B1(\dsmod0.accu1[1] ),
    .X(_03248_));
 sky130_fd_sc_hd__and3_1 _14167_ (.A(\dsmod0.accu1[1] ),
    .B(_03246_),
    .C(_03247_),
    .X(_03249_));
 sky130_fd_sc_hd__a31oi_2 _14168_ (.A1(\dsmod0.accu1[0] ),
    .A2(_03240_),
    .A3(_03248_),
    .B1(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_1 _14169_ (.A(\dsmod0.accu1[2] ),
    .B(_03058_),
    .Y(_03251_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(\dsmod0.accu1[3] ),
    .B(_02963_),
    .Y(_03252_));
 sky130_fd_sc_hd__a211o_1 _14171_ (.A1(_03059_),
    .A2(_03250_),
    .B1(_03251_),
    .C1(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__mux4_1 _14172_ (.A0(_06608_),
    .A1(_06791_),
    .A2(_06917_),
    .A3(_07040_),
    .S0(_07322_),
    .S1(_07315_),
    .X(_03254_));
 sky130_fd_sc_hd__o21a_1 _14173_ (.A1(net32),
    .A2(_03254_),
    .B1(_07168_),
    .X(_03255_));
 sky130_fd_sc_hd__nor2_1 _14174_ (.A(_07314_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__mux2_1 _14175_ (.A0(_02763_),
    .A1(_02573_),
    .S(_06353_),
    .X(_03257_));
 sky130_fd_sc_hd__o21a_1 _14176_ (.A1(_07322_),
    .A2(_02668_),
    .B1(_03053_),
    .X(_03258_));
 sky130_fd_sc_hd__mux4_1 _14177_ (.A0(_02375_),
    .A1(_02374_),
    .A2(_03257_),
    .A3(_03258_),
    .S0(_07315_),
    .S1(_07326_),
    .X(_03259_));
 sky130_fd_sc_hd__a21o_1 _14178_ (.A1(_07314_),
    .A2(_03259_),
    .B1(_07173_),
    .X(_03260_));
 sky130_fd_sc_hd__o221a_2 _14179_ (.A1(_07182_),
    .A2(_03236_),
    .B1(_03256_),
    .B2(_03260_),
    .C1(_07331_),
    .X(_03261_));
 sky130_fd_sc_hd__xnor2_1 _14180_ (.A(\dsmod0.accu1[4] ),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__a21o_1 _14181_ (.A1(_02964_),
    .A2(_03253_),
    .B1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__o21ai_1 _14182_ (.A1(net32),
    .A2(_07319_),
    .B1(_07168_),
    .Y(_03264_));
 sky130_fd_sc_hd__mux4_1 _14183_ (.A0(_02372_),
    .A1(_02375_),
    .A2(_02374_),
    .A3(_03257_),
    .S0(_07165_),
    .S1(_07325_),
    .X(_03265_));
 sky130_fd_sc_hd__mux2_1 _14184_ (.A0(_03264_),
    .A1(_03265_),
    .S(_07170_),
    .X(_03266_));
 sky130_fd_sc_hd__and2_1 _14185_ (.A(_07331_),
    .B(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__nor2_1 _14186_ (.A(\dsmod0.accu1[6] ),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__and3_1 _14187_ (.A(\dsmod0.accu1[6] ),
    .B(_02383_),
    .C(_03266_),
    .X(_03269_));
 sky130_fd_sc_hd__or2_1 _14188_ (.A(_03268_),
    .B(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__mux4_1 _14189_ (.A0(_02174_),
    .A1(_02177_),
    .A2(_02179_),
    .A3(_02574_),
    .S0(_07315_),
    .S1(_07326_),
    .X(_03271_));
 sky130_fd_sc_hd__a21o_1 _14190_ (.A1(_07314_),
    .A2(_03271_),
    .B1(_07328_),
    .X(_03272_));
 sky130_fd_sc_hd__o21a_1 _14191_ (.A1(_07182_),
    .A2(_02573_),
    .B1(_07331_),
    .X(_03273_));
 sky130_fd_sc_hd__and2_1 _14192_ (.A(_03272_),
    .B(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__or2_1 _14193_ (.A(\dsmod0.accu1[7] ),
    .B(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__nand2_1 _14194_ (.A(\dsmod0.accu1[7] ),
    .B(_03274_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _14195_ (.A(_03275_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__a21o_1 _14196_ (.A1(_02383_),
    .A2(_02766_),
    .B1(\dsmod0.accu1[5] ),
    .X(_03278_));
 sky130_fd_sc_hd__and3_1 _14197_ (.A(\dsmod0.accu1[4] ),
    .B(_03278_),
    .C(_03261_),
    .X(_03279_));
 sky130_fd_sc_hd__or2_1 _14198_ (.A(\dsmod0.accu1[6] ),
    .B(_03267_),
    .X(_03280_));
 sky130_fd_sc_hd__o311a_1 _14199_ (.A1(_02769_),
    .A2(_03269_),
    .A3(_03279_),
    .B1(_03275_),
    .C1(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__a21oi_1 _14200_ (.A1(\dsmod0.accu1[7] ),
    .A2(_03274_),
    .B1(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__o41a_1 _14201_ (.A1(_02770_),
    .A2(_03263_),
    .A3(_03270_),
    .A4(_03277_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__or2_1 _14202_ (.A(\dsmod0.accu1[8] ),
    .B(_02378_),
    .X(_03284_));
 sky130_fd_sc_hd__nand2_1 _14203_ (.A(_02379_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__or2_1 _14204_ (.A(\dsmod0.accu1[9] ),
    .B(_02182_),
    .X(_03286_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_02183_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nor4b_1 _14206_ (.A(_03283_),
    .B(_03285_),
    .C(_03287_),
    .D_N(_07334_),
    .Y(_03288_));
 sky130_fd_sc_hd__a21o_1 _14207_ (.A1(\dsmod0.accu1[10] ),
    .A2(_07332_),
    .B1(_07179_),
    .X(_03289_));
 sky130_fd_sc_hd__and2b_1 _14208_ (.A_N(_07178_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a211o_1 _14209_ (.A1(_07334_),
    .A2(_02381_),
    .B1(_03288_),
    .C1(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__a21o_1 _14210_ (.A1(_07314_),
    .A2(_02385_),
    .B1(_07328_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_2 _14211_ (.A1(_07182_),
    .A2(_02371_),
    .B1(_03292_),
    .C1(_02383_),
    .X(_03293_));
 sky130_fd_sc_hd__or2_1 _14212_ (.A(\dsmod0.accu1[13] ),
    .B(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__nand2_1 _14213_ (.A(\dsmod0.accu1[13] ),
    .B(_03293_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _14214_ (.A(_03294_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__inv_2 _14215_ (.A(\dsmod0.accu1[12] ),
    .Y(_03297_));
 sky130_fd_sc_hd__o21a_1 _14216_ (.A1(_06354_),
    .A2(_03255_),
    .B1(_07174_),
    .X(_03298_));
 sky130_fd_sc_hd__a211o_1 _14217_ (.A1(_07173_),
    .A2(_07040_),
    .B1(_03298_),
    .C1(_06356_),
    .X(_03299_));
 sky130_fd_sc_hd__nor2_1 _14218_ (.A(_03297_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__nand2_1 _14219_ (.A(_03297_),
    .B(_03299_),
    .Y(_03301_));
 sky130_fd_sc_hd__or2b_1 _14220_ (.A(_03300_),
    .B_N(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__nor2_1 _14221_ (.A(_03296_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__a21o_1 _14222_ (.A1(\dsmod0.accu1[13] ),
    .A2(_03293_),
    .B1(_03300_),
    .X(_03304_));
 sky130_fd_sc_hd__a22oi_2 _14223_ (.A1(_03291_),
    .A2(_03303_),
    .B1(_03304_),
    .B2(_03294_),
    .Y(_03305_));
 sky130_fd_sc_hd__mux2_1 _14224_ (.A0(_06608_),
    .A1(_06791_),
    .S(_07173_),
    .X(_03306_));
 sky130_fd_sc_hd__nor2_2 _14225_ (.A(_06356_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__and2_1 _14226_ (.A(\dsmod0.accu1[14] ),
    .B(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_1 _14227_ (.A(\dsmod0.accu1[14] ),
    .B(_03307_),
    .Y(_03309_));
 sky130_fd_sc_hd__or2_1 _14228_ (.A(_03308_),
    .B(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_1 _14229_ (.A(_03305_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__inv_2 _14230_ (.A(_06609_),
    .Y(_03312_));
 sky130_fd_sc_hd__o21a_1 _14231_ (.A1(\dsmod0.accu1[15] ),
    .A2(_03312_),
    .B1(_03308_),
    .X(_03313_));
 sky130_fd_sc_hd__a211o_1 _14232_ (.A1(\dsmod0.accu1[15] ),
    .A2(_03312_),
    .B1(_03313_),
    .C1(net18),
    .X(_03314_));
 sky130_fd_sc_hd__a21o_1 _14233_ (.A1(_06610_),
    .A2(_03311_),
    .B1(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__xnor2_1 _14234_ (.A(\dsmod0.mod2_out[1] ),
    .B(\dsmod0.accu3[1] ),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _14235_ (.A(\dsmod0.mod2_out[0] ),
    .B(\dsmod0.accu3[0] ),
    .Y(_03317_));
 sky130_fd_sc_hd__o21ai_1 _14236_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_06348_),
    .Y(_03318_));
 sky130_fd_sc_hd__a21o_1 _14237_ (.A1(\dsmod0.mod2_out[1] ),
    .A2(\dsmod0.accu3[1] ),
    .B1(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__and3_1 _14238_ (.A(_05902_),
    .B(_03315_),
    .C(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _14239_ (.A(_03320_),
    .X(_01986_));
 sky130_fd_sc_hd__clkinv_2 _14240_ (.A(net18),
    .Y(_03321_));
 sky130_fd_sc_hd__buf_4 _14241_ (.A(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__a21o_1 _14242_ (.A1(\dsmod0.mod2_out[0] ),
    .A2(_06349_),
    .B1(\dsmod0.accu3[0] ),
    .X(_03323_));
 sky130_fd_sc_hd__o211a_1 _14243_ (.A1(_03322_),
    .A2(_03317_),
    .B1(_03323_),
    .C1(_05927_),
    .X(_01987_));
 sky130_fd_sc_hd__a21oi_1 _14244_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03318_),
    .Y(_03324_));
 sky130_fd_sc_hd__a21oi_1 _14245_ (.A1(\dsmod0.accu3[1] ),
    .A2(_03322_),
    .B1(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__nor2_1 _14246_ (.A(_05924_),
    .B(_03325_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor3_1 _14247_ (.A(_03321_),
    .B(\dsmod0.mod2_ctr[1] ),
    .C(\dsmod0.mod2_ctr[0] ),
    .Y(_03326_));
 sky130_fd_sc_hd__clkbuf_4 _14248_ (.A(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__buf_2 _14249_ (.A(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__inv_2 _14250_ (.A(\dsmod0.accu1[0] ),
    .Y(_03329_));
 sky130_fd_sc_hd__buf_4 _14251_ (.A(_03327_),
    .X(_03330_));
 sky130_fd_sc_hd__nand2_1 _14252_ (.A(_03329_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__clkbuf_4 _14253_ (.A(_05902_),
    .X(_03332_));
 sky130_fd_sc_hd__o211a_1 _14254_ (.A1(\dsmod0.accu2[0] ),
    .A2(_03328_),
    .B1(_03331_),
    .C1(_03332_),
    .X(_01989_));
 sky130_fd_sc_hd__or3_4 _14255_ (.A(_03321_),
    .B(\dsmod0.mod2_ctr[1] ),
    .C(\dsmod0.mod2_ctr[0] ),
    .X(_03333_));
 sky130_fd_sc_hd__buf_2 _14256_ (.A(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__or2_1 _14257_ (.A(\dsmod0.accu1[1] ),
    .B(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__o211a_1 _14258_ (.A1(\dsmod0.accu2[1] ),
    .A2(_03328_),
    .B1(_03335_),
    .C1(_03332_),
    .X(_01990_));
 sky130_fd_sc_hd__or2_1 _14259_ (.A(\dsmod0.accu1[2] ),
    .B(_03334_),
    .X(_03336_));
 sky130_fd_sc_hd__o211a_1 _14260_ (.A1(\dsmod0.accu2[2] ),
    .A2(_03328_),
    .B1(_03336_),
    .C1(_03332_),
    .X(_01991_));
 sky130_fd_sc_hd__or2_1 _14261_ (.A(\dsmod0.accu1[3] ),
    .B(_03334_),
    .X(_03337_));
 sky130_fd_sc_hd__o211a_1 _14262_ (.A1(\dsmod0.accu2[3] ),
    .A2(_03328_),
    .B1(_03337_),
    .C1(_03332_),
    .X(_01992_));
 sky130_fd_sc_hd__or2_1 _14263_ (.A(\dsmod0.accu1[4] ),
    .B(_03334_),
    .X(_03338_));
 sky130_fd_sc_hd__o211a_1 _14264_ (.A1(\dsmod0.accu2[4] ),
    .A2(_03328_),
    .B1(_03338_),
    .C1(_03332_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _14265_ (.A(_02382_),
    .B(_03330_),
    .Y(_03339_));
 sky130_fd_sc_hd__o211a_1 _14266_ (.A1(\dsmod0.accu2[5] ),
    .A2(_03328_),
    .B1(_03339_),
    .C1(_03332_),
    .X(_01994_));
 sky130_fd_sc_hd__or2_1 _14267_ (.A(\dsmod0.accu1[6] ),
    .B(_03334_),
    .X(_03340_));
 sky130_fd_sc_hd__o211a_1 _14268_ (.A1(\dsmod0.accu2[6] ),
    .A2(_03328_),
    .B1(_03340_),
    .C1(_03332_),
    .X(_01995_));
 sky130_fd_sc_hd__or2_1 _14269_ (.A(\dsmod0.accu1[7] ),
    .B(_03334_),
    .X(_03341_));
 sky130_fd_sc_hd__o211a_1 _14270_ (.A1(\dsmod0.accu2[7] ),
    .A2(_03328_),
    .B1(_03341_),
    .C1(_03332_),
    .X(_01996_));
 sky130_fd_sc_hd__or2_1 _14271_ (.A(\dsmod0.accu1[8] ),
    .B(_03334_),
    .X(_03342_));
 sky130_fd_sc_hd__o211a_1 _14272_ (.A1(\dsmod0.accu2[8] ),
    .A2(_03328_),
    .B1(_03342_),
    .C1(_03332_),
    .X(_01997_));
 sky130_fd_sc_hd__or2_1 _14273_ (.A(\dsmod0.accu1[9] ),
    .B(_03334_),
    .X(_03343_));
 sky130_fd_sc_hd__o211a_1 _14274_ (.A1(\dsmod0.accu2[9] ),
    .A2(_03328_),
    .B1(_03343_),
    .C1(_03332_),
    .X(_01998_));
 sky130_fd_sc_hd__inv_2 _14275_ (.A(\dsmod0.accu1[10] ),
    .Y(_03344_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_03344_),
    .B(_03330_),
    .Y(_03345_));
 sky130_fd_sc_hd__buf_4 _14277_ (.A(_05902_),
    .X(_03346_));
 sky130_fd_sc_hd__o211a_1 _14278_ (.A1(\dsmod0.accu2[10] ),
    .A2(_03330_),
    .B1(_03345_),
    .C1(_03346_),
    .X(_01999_));
 sky130_fd_sc_hd__inv_2 _14279_ (.A(\dsmod0.accu1[11] ),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _14280_ (.A(_03347_),
    .B(_03327_),
    .Y(_03348_));
 sky130_fd_sc_hd__o211a_1 _14281_ (.A1(\dsmod0.accu2[11] ),
    .A2(_03330_),
    .B1(_03348_),
    .C1(_03346_),
    .X(_02000_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_03297_),
    .B(_03327_),
    .Y(_03349_));
 sky130_fd_sc_hd__o211a_1 _14283_ (.A1(\dsmod0.accu2[12] ),
    .A2(_03330_),
    .B1(_03349_),
    .C1(_03346_),
    .X(_02001_));
 sky130_fd_sc_hd__or2_1 _14284_ (.A(\dsmod0.accu1[13] ),
    .B(_03333_),
    .X(_03350_));
 sky130_fd_sc_hd__o211a_1 _14285_ (.A1(\dsmod0.accu2[13] ),
    .A2(_03330_),
    .B1(_03350_),
    .C1(_03346_),
    .X(_02002_));
 sky130_fd_sc_hd__or2_1 _14286_ (.A(\dsmod0.accu1[14] ),
    .B(_03333_),
    .X(_03351_));
 sky130_fd_sc_hd__o211a_1 _14287_ (.A1(\dsmod0.accu2[14] ),
    .A2(_03330_),
    .B1(_03351_),
    .C1(_03346_),
    .X(_02003_));
 sky130_fd_sc_hd__or2_1 _14288_ (.A(\dsmod0.accu1[15] ),
    .B(_03333_),
    .X(_03352_));
 sky130_fd_sc_hd__o211a_1 _14289_ (.A1(\dsmod0.accu2[15] ),
    .A2(_03330_),
    .B1(_03352_),
    .C1(_03346_),
    .X(_02004_));
 sky130_fd_sc_hd__o21ai_1 _14290_ (.A1(\dsmod0.mod2_ctr[1] ),
    .A2(\dsmod0.mod2_ctr[0] ),
    .B1(_06348_),
    .Y(_03353_));
 sky130_fd_sc_hd__buf_4 _14291_ (.A(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__nand2_1 _14292_ (.A(_02383_),
    .B(_03239_),
    .Y(_03355_));
 sky130_fd_sc_hd__mux2_1 _14293_ (.A0(\dsmod0.accu1[0] ),
    .A1(\dsmod0.accu2[0] ),
    .S(_06348_),
    .X(_03356_));
 sky130_fd_sc_hd__o21a_1 _14294_ (.A1(\dsmod0.mod2_ctr[1] ),
    .A2(\dsmod0.mod2_ctr[0] ),
    .B1(net18),
    .X(_03357_));
 sky130_fd_sc_hd__buf_4 _14295_ (.A(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__a21o_1 _14296_ (.A1(_03355_),
    .A2(_03356_),
    .B1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__nor2_1 _14297_ (.A(_03355_),
    .B(_03356_),
    .Y(_03360_));
 sky130_fd_sc_hd__buf_4 _14298_ (.A(_05902_),
    .X(_03361_));
 sky130_fd_sc_hd__o221a_1 _14299_ (.A1(\dsmod0.accu1[0] ),
    .A2(_03354_),
    .B1(_03359_),
    .B2(_03360_),
    .C1(_03361_),
    .X(_02005_));
 sky130_fd_sc_hd__and2_1 _14300_ (.A(\dsmod0.accu1[1] ),
    .B(_03358_),
    .X(_03362_));
 sky130_fd_sc_hd__inv_2 _14301_ (.A(\dsmod0.accu2[1] ),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3_1 _14302_ (.A(\dsmod0.accu1[0] ),
    .B(_03246_),
    .C(_03247_),
    .Y(_03364_));
 sky130_fd_sc_hd__a21o_1 _14303_ (.A1(_03246_),
    .A2(_03247_),
    .B1(\dsmod0.accu1[0] ),
    .X(_03365_));
 sky130_fd_sc_hd__and3_1 _14304_ (.A(_03363_),
    .B(_03364_),
    .C(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_1 _14305_ (.A1(_03364_),
    .A2(_03365_),
    .B1(_03363_),
    .Y(_03367_));
 sky130_fd_sc_hd__nor2_1 _14306_ (.A(_03366_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _14307_ (.A(\dsmod0.accu2[0] ),
    .B(_03355_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(_03368_),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__or2_1 _14309_ (.A(_03368_),
    .B(_03369_),
    .X(_03371_));
 sky130_fd_sc_hd__nor2_1 _14310_ (.A(_03329_),
    .B(_03355_),
    .Y(_03372_));
 sky130_fd_sc_hd__or2b_1 _14311_ (.A(_03249_),
    .B_N(_03248_),
    .X(_03373_));
 sky130_fd_sc_hd__xnor2_1 _14312_ (.A(_03372_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__a32o_1 _14313_ (.A1(_03327_),
    .A2(_03370_),
    .A3(_03371_),
    .B1(_03374_),
    .B2(_03322_),
    .X(_03375_));
 sky130_fd_sc_hd__o21a_1 _14314_ (.A1(_03362_),
    .A2(_03375_),
    .B1(_05927_),
    .X(_02006_));
 sky130_fd_sc_hd__o21ba_1 _14315_ (.A1(_06356_),
    .A2(_03057_),
    .B1_N(\dsmod0.accu1[1] ),
    .X(_03376_));
 sky130_fd_sc_hd__and3b_1 _14316_ (.A_N(_03057_),
    .B(\dsmod0.accu1[1] ),
    .C(_07331_),
    .X(_03377_));
 sky130_fd_sc_hd__or3_1 _14317_ (.A(\dsmod0.accu2[2] ),
    .B(_03376_),
    .C(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__o21ai_1 _14318_ (.A1(_03376_),
    .A2(_03377_),
    .B1(\dsmod0.accu2[2] ),
    .Y(_03379_));
 sky130_fd_sc_hd__a21bo_1 _14319_ (.A1(_03363_),
    .A2(_03365_),
    .B1_N(_03364_),
    .X(_03380_));
 sky130_fd_sc_hd__and3_1 _14320_ (.A(_03378_),
    .B(_03379_),
    .C(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__a21oi_1 _14321_ (.A1(_03378_),
    .A2(_03379_),
    .B1(_03380_),
    .Y(_03382_));
 sky130_fd_sc_hd__or3_1 _14322_ (.A(_03370_),
    .B(_03381_),
    .C(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__o21ai_1 _14323_ (.A1(_03381_),
    .A2(_03382_),
    .B1(_03370_),
    .Y(_03384_));
 sky130_fd_sc_hd__and2_1 _14324_ (.A(\dsmod0.accu1[2] ),
    .B(_03058_),
    .X(_03385_));
 sky130_fd_sc_hd__o21ai_1 _14325_ (.A1(_03385_),
    .A2(_03251_),
    .B1(_03250_),
    .Y(_03386_));
 sky130_fd_sc_hd__or3_1 _14326_ (.A(_03385_),
    .B(_03251_),
    .C(_03250_),
    .X(_03387_));
 sky130_fd_sc_hd__a31o_1 _14327_ (.A1(_03321_),
    .A2(_03386_),
    .A3(_03387_),
    .B1(_03357_),
    .X(_03388_));
 sky130_fd_sc_hd__a31o_1 _14328_ (.A1(_06349_),
    .A2(_03383_),
    .A3(_03384_),
    .B1(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__o211a_1 _14329_ (.A1(\dsmod0.accu1[2] ),
    .A2(_03354_),
    .B1(_03389_),
    .C1(_03346_),
    .X(_02007_));
 sky130_fd_sc_hd__a21o_1 _14330_ (.A1(_03378_),
    .A2(_03379_),
    .B1(_03380_),
    .X(_03390_));
 sky130_fd_sc_hd__a31oi_2 _14331_ (.A1(_03368_),
    .A2(_03369_),
    .A3(_03390_),
    .B1(_03381_),
    .Y(_03391_));
 sky130_fd_sc_hd__nor3_1 _14332_ (.A(\dsmod0.accu2[2] ),
    .B(_03376_),
    .C(_03377_),
    .Y(_03392_));
 sky130_fd_sc_hd__xnor2_1 _14333_ (.A(\dsmod0.accu1[2] ),
    .B(_02963_),
    .Y(_03393_));
 sky130_fd_sc_hd__xor2_1 _14334_ (.A(\dsmod0.accu2[3] ),
    .B(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__nor3_1 _14335_ (.A(_03377_),
    .B(_03392_),
    .C(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__o21a_1 _14336_ (.A1(_03377_),
    .A2(_03392_),
    .B1(_03394_),
    .X(_03396_));
 sky130_fd_sc_hd__nor2_1 _14337_ (.A(_03395_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__xnor2_1 _14338_ (.A(_03391_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__inv_2 _14339_ (.A(_03252_),
    .Y(_03399_));
 sky130_fd_sc_hd__a21o_1 _14340_ (.A1(_03059_),
    .A2(_03250_),
    .B1(_03251_),
    .X(_03400_));
 sky130_fd_sc_hd__a21oi_1 _14341_ (.A1(_02964_),
    .A2(_03399_),
    .B1(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__and3_1 _14342_ (.A(_02964_),
    .B(_03399_),
    .C(_03400_),
    .X(_03402_));
 sky130_fd_sc_hd__or3_1 _14343_ (.A(_06348_),
    .B(_03401_),
    .C(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__a22o_1 _14344_ (.A1(_06349_),
    .A2(_03398_),
    .B1(_03403_),
    .B2(_03334_),
    .X(_03404_));
 sky130_fd_sc_hd__o211a_1 _14345_ (.A1(\dsmod0.accu1[3] ),
    .A2(_03354_),
    .B1(_03404_),
    .C1(_03346_),
    .X(_02008_));
 sky130_fd_sc_hd__xnor2_1 _14346_ (.A(\dsmod0.accu1[3] ),
    .B(_03261_),
    .Y(_03405_));
 sky130_fd_sc_hd__xor2_1 _14347_ (.A(\dsmod0.accu2[4] ),
    .B(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__and3_1 _14348_ (.A(\dsmod0.accu1[2] ),
    .B(_02383_),
    .C(_02962_),
    .X(_03407_));
 sky130_fd_sc_hd__o21bai_1 _14349_ (.A1(\dsmod0.accu2[3] ),
    .A2(_03393_),
    .B1_N(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__xor2_1 _14350_ (.A(_03406_),
    .B(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__inv_2 _14351_ (.A(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ba_2 _14352_ (.A1(_03395_),
    .A2(_03391_),
    .B1_N(_03396_),
    .X(_03411_));
 sky130_fd_sc_hd__nand2_1 _14353_ (.A(_03410_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__or2_1 _14354_ (.A(_03410_),
    .B(_03411_),
    .X(_03413_));
 sky130_fd_sc_hd__and3_1 _14355_ (.A(_03327_),
    .B(_03412_),
    .C(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__nand3_1 _14356_ (.A(_02964_),
    .B(_03253_),
    .C(_03262_),
    .Y(_03415_));
 sky130_fd_sc_hd__a32o_1 _14357_ (.A1(_03322_),
    .A2(_03263_),
    .A3(_03415_),
    .B1(_03358_),
    .B2(\dsmod0.accu1[4] ),
    .X(_03416_));
 sky130_fd_sc_hd__o21a_1 _14358_ (.A1(_03414_),
    .A2(_03416_),
    .B1(_05927_),
    .X(_02009_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_03406_),
    .B(_03408_),
    .Y(_03417_));
 sky130_fd_sc_hd__and2_1 _14360_ (.A(\dsmod0.accu1[3] ),
    .B(_03261_),
    .X(_03418_));
 sky130_fd_sc_hd__nor2_1 _14361_ (.A(\dsmod0.accu2[4] ),
    .B(_03405_),
    .Y(_03419_));
 sky130_fd_sc_hd__a21oi_1 _14362_ (.A1(_02383_),
    .A2(_02766_),
    .B1(\dsmod0.accu1[4] ),
    .Y(_03420_));
 sky130_fd_sc_hd__and3_1 _14363_ (.A(\dsmod0.accu1[4] ),
    .B(_02383_),
    .C(_02766_),
    .X(_03421_));
 sky130_fd_sc_hd__nor2_1 _14364_ (.A(_03420_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__xnor2_1 _14365_ (.A(\dsmod0.accu2[5] ),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__o21ai_2 _14366_ (.A1(_03418_),
    .A2(_03419_),
    .B1(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor3_2 _14368_ (.A(_03418_),
    .B(_03419_),
    .C(_03423_),
    .Y(_03426_));
 sky130_fd_sc_hd__a211o_1 _14369_ (.A1(_03417_),
    .A2(_03413_),
    .B1(_03425_),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__o211a_1 _14370_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03417_),
    .C1(_03413_),
    .X(_03428_));
 sky130_fd_sc_hd__nor2_1 _14371_ (.A(_03322_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__a21bo_1 _14372_ (.A1(\dsmod0.accu1[4] ),
    .A2(_03261_),
    .B1_N(_03263_),
    .X(_03430_));
 sky130_fd_sc_hd__xnor2_1 _14373_ (.A(_02770_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__a221o_1 _14374_ (.A1(_03427_),
    .A2(_03429_),
    .B1(_03431_),
    .B2(_03322_),
    .C1(_03358_),
    .X(_03432_));
 sky130_fd_sc_hd__o211a_1 _14375_ (.A1(\dsmod0.accu1[5] ),
    .A2(_03354_),
    .B1(_03432_),
    .C1(_03346_),
    .X(_02010_));
 sky130_fd_sc_hd__xnor2_1 _14376_ (.A(_02382_),
    .B(_03267_),
    .Y(_03433_));
 sky130_fd_sc_hd__xnor2_1 _14377_ (.A(\dsmod0.accu2[6] ),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__inv_2 _14378_ (.A(\dsmod0.accu2[5] ),
    .Y(_03435_));
 sky130_fd_sc_hd__a21o_1 _14379_ (.A1(_03435_),
    .A2(_03422_),
    .B1(_03421_),
    .X(_03436_));
 sky130_fd_sc_hd__xnor2_1 _14380_ (.A(_03434_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__nand3b_2 _14381_ (.A_N(_03426_),
    .B(_03409_),
    .C(_03424_),
    .Y(_03438_));
 sky130_fd_sc_hd__a21o_1 _14382_ (.A1(_03417_),
    .A2(_03424_),
    .B1(_03426_),
    .X(_03439_));
 sky130_fd_sc_hd__o21a_1 _14383_ (.A1(_03411_),
    .A2(_03438_),
    .B1(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__or2_1 _14384_ (.A(_03437_),
    .B(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__nand2_1 _14385_ (.A(_03437_),
    .B(_03440_),
    .Y(_03442_));
 sky130_fd_sc_hd__and3_1 _14386_ (.A(_03327_),
    .B(_03441_),
    .C(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__nor2_1 _14387_ (.A(_02770_),
    .B(_03263_),
    .Y(_03444_));
 sky130_fd_sc_hd__or3_1 _14388_ (.A(_02769_),
    .B(_03444_),
    .C(_03279_),
    .X(_03445_));
 sky130_fd_sc_hd__xnor2_1 _14389_ (.A(_03270_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__a22o_1 _14390_ (.A1(\dsmod0.accu1[6] ),
    .A2(_03358_),
    .B1(_03446_),
    .B2(_03322_),
    .X(_03447_));
 sky130_fd_sc_hd__o21a_1 _14391_ (.A1(_03443_),
    .A2(_03447_),
    .B1(_05927_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_1 _14392_ (.A(_03434_),
    .B(_03436_),
    .Y(_03448_));
 sky130_fd_sc_hd__inv_2 _14393_ (.A(\dsmod0.accu2[6] ),
    .Y(_03449_));
 sky130_fd_sc_hd__and3_1 _14394_ (.A(\dsmod0.accu1[5] ),
    .B(_02383_),
    .C(_03266_),
    .X(_03450_));
 sky130_fd_sc_hd__a21o_1 _14395_ (.A1(_03449_),
    .A2(_03433_),
    .B1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_2 _14396_ (.A(\dsmod0.accu1[6] ),
    .B(_03274_),
    .Y(_03452_));
 sky130_fd_sc_hd__xor2_2 _14397_ (.A(\dsmod0.accu2[7] ),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__xnor2_1 _14398_ (.A(_03451_),
    .B(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21oi_1 _14399_ (.A1(_03448_),
    .A2(_03441_),
    .B1(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__a31o_1 _14400_ (.A1(_03448_),
    .A2(_03441_),
    .A3(_03454_),
    .B1(_03321_),
    .X(_03456_));
 sky130_fd_sc_hd__a21oi_1 _14401_ (.A1(_03280_),
    .A2(_03445_),
    .B1(_03269_),
    .Y(_03457_));
 sky130_fd_sc_hd__xnor2_1 _14402_ (.A(_03277_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__o221ai_1 _14403_ (.A1(_03455_),
    .A2(_03456_),
    .B1(_03458_),
    .B2(_06349_),
    .C1(_03354_),
    .Y(_03459_));
 sky130_fd_sc_hd__o211a_1 _14404_ (.A1(\dsmod0.accu1[7] ),
    .A2(_03354_),
    .B1(_03459_),
    .C1(_03346_),
    .X(_02012_));
 sky130_fd_sc_hd__or2_1 _14405_ (.A(_03283_),
    .B(_03285_),
    .X(_03460_));
 sky130_fd_sc_hd__nand2_1 _14406_ (.A(_03322_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_1 _14407_ (.A1(_03283_),
    .A2(_03285_),
    .B1(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__or2_1 _14408_ (.A(_03437_),
    .B(_03454_),
    .X(_03463_));
 sky130_fd_sc_hd__a2111o_1 _14409_ (.A1(_03417_),
    .A2(_03424_),
    .B1(_03426_),
    .C1(_03437_),
    .D1(_03454_),
    .X(_03464_));
 sky130_fd_sc_hd__a22o_1 _14410_ (.A1(_03434_),
    .A2(_03436_),
    .B1(_03451_),
    .B2(_03453_),
    .X(_03465_));
 sky130_fd_sc_hd__o21ai_1 _14411_ (.A1(_03451_),
    .A2(_03453_),
    .B1(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__o311ai_4 _14412_ (.A1(_03411_),
    .A2(_03438_),
    .A3(_03463_),
    .B1(_03464_),
    .C1(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__and3_1 _14413_ (.A(\dsmod0.accu1[6] ),
    .B(_03272_),
    .C(_03273_),
    .X(_03468_));
 sky130_fd_sc_hd__nor2_1 _14414_ (.A(\dsmod0.accu2[7] ),
    .B(_03452_),
    .Y(_03469_));
 sky130_fd_sc_hd__xnor2_1 _14415_ (.A(\dsmod0.accu1[7] ),
    .B(_02378_),
    .Y(_03470_));
 sky130_fd_sc_hd__xor2_1 _14416_ (.A(\dsmod0.accu2[8] ),
    .B(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__o21ai_1 _14417_ (.A1(_03468_),
    .A2(_03469_),
    .B1(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__or3_1 _14418_ (.A(_03468_),
    .B(_03469_),
    .C(_03471_),
    .X(_03473_));
 sky130_fd_sc_hd__and2_1 _14419_ (.A(_03472_),
    .B(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__or2_1 _14420_ (.A(_03467_),
    .B(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_03467_),
    .B(_03474_),
    .Y(_03476_));
 sky130_fd_sc_hd__a32o_1 _14422_ (.A1(_03327_),
    .A2(_03475_),
    .A3(_03476_),
    .B1(_03358_),
    .B2(\dsmod0.accu1[8] ),
    .X(_03477_));
 sky130_fd_sc_hd__o21a_1 _14423_ (.A1(_03462_),
    .A2(_03477_),
    .B1(_05927_),
    .X(_02013_));
 sky130_fd_sc_hd__and2_1 _14424_ (.A(\dsmod0.accu1[7] ),
    .B(_02378_),
    .X(_03478_));
 sky130_fd_sc_hd__nor2_1 _14425_ (.A(\dsmod0.accu2[8] ),
    .B(_03470_),
    .Y(_03479_));
 sky130_fd_sc_hd__xnor2_1 _14426_ (.A(\dsmod0.accu1[8] ),
    .B(_02182_),
    .Y(_03480_));
 sky130_fd_sc_hd__xor2_1 _14427_ (.A(\dsmod0.accu2[9] ),
    .B(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__o21ai_1 _14428_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__or3_1 _14429_ (.A(_03478_),
    .B(_03479_),
    .C(_03481_),
    .X(_03483_));
 sky130_fd_sc_hd__and2_1 _14430_ (.A(_03482_),
    .B(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__a21bo_1 _14431_ (.A1(_03467_),
    .A2(_03474_),
    .B1_N(_03472_),
    .X(_03485_));
 sky130_fd_sc_hd__o21ai_1 _14432_ (.A1(_03484_),
    .A2(_03485_),
    .B1(_06349_),
    .Y(_03486_));
 sky130_fd_sc_hd__a21oi_1 _14433_ (.A1(_03484_),
    .A2(_03485_),
    .B1(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__nand2_1 _14434_ (.A(_02379_),
    .B(_03460_),
    .Y(_03488_));
 sky130_fd_sc_hd__xor2_1 _14435_ (.A(_03488_),
    .B(_03287_),
    .X(_03489_));
 sky130_fd_sc_hd__a21oi_1 _14436_ (.A1(_03322_),
    .A2(_03489_),
    .B1(_03327_),
    .Y(_03490_));
 sky130_fd_sc_hd__o221a_1 _14437_ (.A1(\dsmod0.accu1[9] ),
    .A2(_03354_),
    .B1(_03487_),
    .B2(_03490_),
    .C1(_03361_),
    .X(_02014_));
 sky130_fd_sc_hd__a21o_1 _14438_ (.A1(_02379_),
    .A2(_03460_),
    .B1(_02380_),
    .X(_03491_));
 sky130_fd_sc_hd__and3_1 _14439_ (.A(_07333_),
    .B(_02183_),
    .C(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__a21oi_1 _14440_ (.A1(_02183_),
    .A2(_03491_),
    .B1(_07333_),
    .Y(_03493_));
 sky130_fd_sc_hd__or3_1 _14441_ (.A(_06348_),
    .B(_03492_),
    .C(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__xor2_1 _14442_ (.A(\dsmod0.accu1[9] ),
    .B(_07332_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _14443_ (.A(\dsmod0.accu2[10] ),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand2_1 _14444_ (.A(\dsmod0.accu1[8] ),
    .B(_02182_),
    .Y(_03497_));
 sky130_fd_sc_hd__o21ai_1 _14445_ (.A1(\dsmod0.accu2[9] ),
    .A2(_03480_),
    .B1(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__xor2_1 _14446_ (.A(_03496_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__and2_1 _14447_ (.A(_03474_),
    .B(_03484_),
    .X(_03500_));
 sky130_fd_sc_hd__a21boi_1 _14448_ (.A1(_03472_),
    .A2(_03482_),
    .B1_N(_03483_),
    .Y(_03501_));
 sky130_fd_sc_hd__a21o_1 _14449_ (.A1(_03467_),
    .A2(_03500_),
    .B1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__and2_1 _14450_ (.A(_03499_),
    .B(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__nor2_1 _14451_ (.A(_03499_),
    .B(_03502_),
    .Y(_03504_));
 sky130_fd_sc_hd__o32a_1 _14452_ (.A1(_03333_),
    .A2(_03503_),
    .A3(_03504_),
    .B1(_03353_),
    .B2(_03344_),
    .X(_03505_));
 sky130_fd_sc_hd__a21oi_1 _14453_ (.A1(_03494_),
    .A2(_03505_),
    .B1(_05924_),
    .Y(_02015_));
 sky130_fd_sc_hd__and2_1 _14454_ (.A(_03496_),
    .B(_03498_),
    .X(_03506_));
 sky130_fd_sc_hd__inv_2 _14455_ (.A(\dsmod0.accu2[10] ),
    .Y(_03507_));
 sky130_fd_sc_hd__and2_1 _14456_ (.A(\dsmod0.accu1[9] ),
    .B(_07332_),
    .X(_03508_));
 sky130_fd_sc_hd__a21o_1 _14457_ (.A1(_03507_),
    .A2(_03495_),
    .B1(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__xnor2_1 _14458_ (.A(\dsmod0.accu1[10] ),
    .B(_07177_),
    .Y(_03510_));
 sky130_fd_sc_hd__xor2_2 _14459_ (.A(\dsmod0.accu2[11] ),
    .B(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__xor2_1 _14460_ (.A(_03509_),
    .B(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__o21ai_1 _14461_ (.A1(_03506_),
    .A2(_03503_),
    .B1(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__o31a_1 _14462_ (.A1(_03506_),
    .A2(_03503_),
    .A3(_03512_),
    .B1(_06348_),
    .X(_03514_));
 sky130_fd_sc_hd__a21o_1 _14463_ (.A1(\dsmod0.accu1[10] ),
    .A2(_07332_),
    .B1(_03493_),
    .X(_03515_));
 sky130_fd_sc_hd__xnor2_1 _14464_ (.A(_07180_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__a221o_1 _14465_ (.A1(_03513_),
    .A2(_03514_),
    .B1(_03516_),
    .B2(_03322_),
    .C1(_03358_),
    .X(_03517_));
 sky130_fd_sc_hd__o211a_1 _14466_ (.A1(\dsmod0.accu1[11] ),
    .A2(_03354_),
    .B1(_03517_),
    .C1(_03361_),
    .X(_02016_));
 sky130_fd_sc_hd__inv_2 _14467_ (.A(_03302_),
    .Y(_03518_));
 sky130_fd_sc_hd__a21oi_1 _14468_ (.A1(_03291_),
    .A2(_03518_),
    .B1(_06348_),
    .Y(_03519_));
 sky130_fd_sc_hd__o21a_1 _14469_ (.A1(_03291_),
    .A2(_03518_),
    .B1(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__and3_1 _14470_ (.A(\dsmod0.accu1[10] ),
    .B(_07175_),
    .C(_07176_),
    .X(_03521_));
 sky130_fd_sc_hd__nor2_1 _14471_ (.A(\dsmod0.accu2[11] ),
    .B(_03510_),
    .Y(_03522_));
 sky130_fd_sc_hd__nor2_1 _14472_ (.A(_03347_),
    .B(_03299_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _14473_ (.A(_03347_),
    .B(_03299_),
    .Y(_03524_));
 sky130_fd_sc_hd__or2b_1 _14474_ (.A(_03523_),
    .B_N(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__nor2_1 _14475_ (.A(\dsmod0.accu2[12] ),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__and2_1 _14476_ (.A(\dsmod0.accu2[12] ),
    .B(_03525_),
    .X(_03527_));
 sky130_fd_sc_hd__nor2_1 _14477_ (.A(_03526_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21a_1 _14478_ (.A1(_03521_),
    .A2(_03522_),
    .B1(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__nor3_1 _14479_ (.A(_03521_),
    .B(_03522_),
    .C(_03528_),
    .Y(_03530_));
 sky130_fd_sc_hd__nor2_1 _14480_ (.A(_03529_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__and2_1 _14481_ (.A(_03499_),
    .B(_03512_),
    .X(_03532_));
 sky130_fd_sc_hd__o21a_1 _14482_ (.A1(_03509_),
    .A2(_03511_),
    .B1(_03506_),
    .X(_03533_));
 sky130_fd_sc_hd__a221o_1 _14483_ (.A1(_03509_),
    .A2(_03511_),
    .B1(_03532_),
    .B2(_03501_),
    .C1(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__a31o_1 _14484_ (.A1(_03467_),
    .A2(_03500_),
    .A3(_03532_),
    .B1(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__and2_1 _14485_ (.A(_03531_),
    .B(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__o21ai_1 _14486_ (.A1(_03531_),
    .A2(_03535_),
    .B1(_03326_),
    .Y(_03537_));
 sky130_fd_sc_hd__a2bb2o_1 _14487_ (.A1_N(_03536_),
    .A2_N(_03537_),
    .B1(\dsmod0.accu1[12] ),
    .B2(_03358_),
    .X(_03538_));
 sky130_fd_sc_hd__o21a_1 _14488_ (.A1(_03520_),
    .A2(_03538_),
    .B1(_05927_),
    .X(_02017_));
 sky130_fd_sc_hd__a21oi_1 _14489_ (.A1(_03291_),
    .A2(_03518_),
    .B1(_03300_),
    .Y(_03539_));
 sky130_fd_sc_hd__xor2_1 _14490_ (.A(_03296_),
    .B(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__nor2_1 _14491_ (.A(\dsmod0.accu1[12] ),
    .B(_03293_),
    .Y(_03541_));
 sky130_fd_sc_hd__and2_1 _14492_ (.A(\dsmod0.accu1[12] ),
    .B(_03293_),
    .X(_03542_));
 sky130_fd_sc_hd__or2_1 _14493_ (.A(_03541_),
    .B(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__nor2_1 _14494_ (.A(\dsmod0.accu2[13] ),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__and2_1 _14495_ (.A(\dsmod0.accu2[13] ),
    .B(_03543_),
    .X(_03545_));
 sky130_fd_sc_hd__nor2_1 _14496_ (.A(_03544_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__o21a_1 _14497_ (.A1(_03523_),
    .A2(_03526_),
    .B1(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__or3_1 _14498_ (.A(_03523_),
    .B(_03526_),
    .C(_03546_),
    .X(_03548_));
 sky130_fd_sc_hd__and2b_1 _14499_ (.A_N(_03547_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__nor2_1 _14500_ (.A(_03529_),
    .B(_03536_),
    .Y(_03550_));
 sky130_fd_sc_hd__and2_1 _14501_ (.A(_03549_),
    .B(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__o21ai_1 _14502_ (.A1(_03549_),
    .A2(_03550_),
    .B1(_03327_),
    .Y(_03552_));
 sky130_fd_sc_hd__o221a_1 _14503_ (.A1(\dsmod0.accu1[13] ),
    .A2(_03354_),
    .B1(_03551_),
    .B2(_03552_),
    .C1(_05902_),
    .X(_03553_));
 sky130_fd_sc_hd__o21a_1 _14504_ (.A1(_06349_),
    .A2(_03540_),
    .B1(_03553_),
    .X(_02018_));
 sky130_fd_sc_hd__nand2_1 _14505_ (.A(_03305_),
    .B(_03310_),
    .Y(_03554_));
 sky130_fd_sc_hd__or3b_1 _14506_ (.A(_06348_),
    .B(_03311_),
    .C_N(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__and2_1 _14507_ (.A(\dsmod0.accu1[13] ),
    .B(_03307_),
    .X(_03556_));
 sky130_fd_sc_hd__nor2_1 _14508_ (.A(\dsmod0.accu1[13] ),
    .B(_03307_),
    .Y(_03557_));
 sky130_fd_sc_hd__or2_1 _14509_ (.A(_03556_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_1 _14510_ (.A(\dsmod0.accu2[14] ),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__and2_1 _14511_ (.A(\dsmod0.accu2[14] ),
    .B(_03558_),
    .X(_03560_));
 sky130_fd_sc_hd__nor2_1 _14512_ (.A(_03559_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__o21a_1 _14513_ (.A1(_03542_),
    .A2(_03544_),
    .B1(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__or3_1 _14514_ (.A(_03542_),
    .B(_03544_),
    .C(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__and2b_1 _14515_ (.A_N(_03562_),
    .B(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__o21a_1 _14516_ (.A1(_03529_),
    .A2(_03547_),
    .B1(_03548_),
    .X(_03565_));
 sky130_fd_sc_hd__a31o_1 _14517_ (.A1(_03531_),
    .A2(_03535_),
    .A3(_03549_),
    .B1(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__xnor2_1 _14518_ (.A(_03564_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__o2bb2a_1 _14519_ (.A1_N(\dsmod0.accu1[14] ),
    .A2_N(_03358_),
    .B1(_03567_),
    .B2(_03333_),
    .X(_03568_));
 sky130_fd_sc_hd__a21oi_1 _14520_ (.A1(_03555_),
    .A2(_03568_),
    .B1(_05924_),
    .Y(_02019_));
 sky130_fd_sc_hd__o21ai_1 _14521_ (.A1(_03308_),
    .A2(_03311_),
    .B1(_06610_),
    .Y(_03569_));
 sky130_fd_sc_hd__o31a_1 _14522_ (.A1(_06610_),
    .A2(_03308_),
    .A3(_03311_),
    .B1(_03321_),
    .X(_03570_));
 sky130_fd_sc_hd__a21oi_1 _14523_ (.A1(_03563_),
    .A2(_03566_),
    .B1(_03562_),
    .Y(_03571_));
 sky130_fd_sc_hd__xnor2_1 _14524_ (.A(\dsmod0.accu1[14] ),
    .B(_06609_),
    .Y(_03572_));
 sky130_fd_sc_hd__and2b_1 _14525_ (.A_N(\dsmod0.accu2[15] ),
    .B(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__and2b_1 _14526_ (.A_N(_03572_),
    .B(\dsmod0.accu2[15] ),
    .X(_03574_));
 sky130_fd_sc_hd__nor2_1 _14527_ (.A(_03573_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__nor3_1 _14528_ (.A(_03556_),
    .B(_03559_),
    .C(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__o21a_1 _14529_ (.A1(_03556_),
    .A2(_03559_),
    .B1(_03575_),
    .X(_03577_));
 sky130_fd_sc_hd__nor2_1 _14530_ (.A(_03576_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__xnor2_1 _14531_ (.A(_03571_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__a221o_1 _14532_ (.A1(_03569_),
    .A2(_03570_),
    .B1(_03579_),
    .B2(_06348_),
    .C1(_03358_),
    .X(_03580_));
 sky130_fd_sc_hd__o211a_1 _14533_ (.A1(\dsmod0.accu1[15] ),
    .A2(_03354_),
    .B1(_03580_),
    .C1(_03361_),
    .X(_02020_));
 sky130_fd_sc_hd__nor2_8 _14534_ (.A(_03919_),
    .B(_05588_),
    .Y(_03581_));
 sky130_fd_sc_hd__buf_6 _14535_ (.A(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__mux2_1 _14536_ (.A0(\fifo0.fifo_store[39][0] ),
    .A1(_06283_),
    .S(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_1 _14537_ (.A(_03583_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _14538_ (.A0(\fifo0.fifo_store[39][1] ),
    .A1(_06287_),
    .S(_03582_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _14539_ (.A(_03584_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _14540_ (.A0(\fifo0.fifo_store[39][2] ),
    .A1(_06310_),
    .S(_03582_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _14541_ (.A(_03585_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _14542_ (.A0(\fifo0.fifo_store[39][3] ),
    .A1(_06312_),
    .S(_03582_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _14543_ (.A(_03586_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _14544_ (.A0(\fifo0.fifo_store[39][4] ),
    .A1(_06314_),
    .S(_03582_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _14545_ (.A(_03587_),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _14546_ (.A0(\fifo0.fifo_store[39][5] ),
    .A1(_03884_),
    .S(_03582_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _14547_ (.A(_03588_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _14548_ (.A0(\fifo0.fifo_store[39][6] ),
    .A1(_06317_),
    .S(_03582_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _14549_ (.A(_03589_),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _14550_ (.A0(\fifo0.fifo_store[39][7] ),
    .A1(_03890_),
    .S(_03582_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _14551_ (.A(_03590_),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _14552_ (.A0(\fifo0.fifo_store[39][8] ),
    .A1(_06320_),
    .S(_03582_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _14553_ (.A(_03591_),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _14554_ (.A0(\fifo0.fifo_store[39][9] ),
    .A1(_06322_),
    .S(_03582_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _14555_ (.A(_03592_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _14556_ (.A0(\fifo0.fifo_store[39][10] ),
    .A1(_03899_),
    .S(_03581_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _14557_ (.A(_03593_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _14558_ (.A0(\fifo0.fifo_store[39][11] ),
    .A1(_03902_),
    .S(_03581_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _14559_ (.A(_03594_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _14560_ (.A0(\fifo0.fifo_store[39][12] ),
    .A1(_06278_),
    .S(_03581_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _14561_ (.A(_03595_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _14562_ (.A0(\fifo0.fifo_store[39][13] ),
    .A1(_06300_),
    .S(_03581_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _14563_ (.A(_03596_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _14564_ (.A0(\fifo0.fifo_store[39][14] ),
    .A1(_06302_),
    .S(_03581_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _14565_ (.A(_03597_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _14566_ (.A0(\fifo0.fifo_store[39][15] ),
    .A1(_06304_),
    .S(_03581_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _14567_ (.A(_03598_),
    .X(_02036_));
 sky130_fd_sc_hd__nor2_8 _14568_ (.A(_03919_),
    .B(_04317_),
    .Y(_03599_));
 sky130_fd_sc_hd__buf_8 _14569_ (.A(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__mux2_1 _14570_ (.A0(\fifo0.fifo_store[119][0] ),
    .A1(_06283_),
    .S(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _14571_ (.A(_03601_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _14572_ (.A0(\fifo0.fifo_store[119][1] ),
    .A1(_06287_),
    .S(_03600_),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _14573_ (.A(_03602_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _14574_ (.A0(\fifo0.fifo_store[119][2] ),
    .A1(_06310_),
    .S(_03600_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _14575_ (.A(_03603_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _14576_ (.A0(\fifo0.fifo_store[119][3] ),
    .A1(_06312_),
    .S(_03600_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_1 _14577_ (.A(_03604_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\fifo0.fifo_store[119][4] ),
    .A1(_06314_),
    .S(_03600_),
    .X(_03605_));
 sky130_fd_sc_hd__clkbuf_1 _14579_ (.A(_03605_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _14580_ (.A0(\fifo0.fifo_store[119][5] ),
    .A1(_03884_),
    .S(_03600_),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_1 _14581_ (.A(_03606_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _14582_ (.A0(\fifo0.fifo_store[119][6] ),
    .A1(_06317_),
    .S(_03600_),
    .X(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _14583_ (.A(_03607_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _14584_ (.A0(\fifo0.fifo_store[119][7] ),
    .A1(_03890_),
    .S(_03600_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _14585_ (.A(_03608_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _14586_ (.A0(\fifo0.fifo_store[119][8] ),
    .A1(_06320_),
    .S(_03600_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _14587_ (.A(_03609_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _14588_ (.A0(\fifo0.fifo_store[119][9] ),
    .A1(_06322_),
    .S(_03600_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _14589_ (.A(_03610_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _14590_ (.A0(\fifo0.fifo_store[119][10] ),
    .A1(_03899_),
    .S(_03599_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _14591_ (.A(_03611_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _14592_ (.A0(\fifo0.fifo_store[119][11] ),
    .A1(_03902_),
    .S(_03599_),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _14593_ (.A(_03612_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _14594_ (.A0(\fifo0.fifo_store[119][12] ),
    .A1(_06278_),
    .S(_03599_),
    .X(_03613_));
 sky130_fd_sc_hd__clkbuf_1 _14595_ (.A(_03613_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _14596_ (.A0(\fifo0.fifo_store[119][13] ),
    .A1(_06300_),
    .S(_03599_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _14597_ (.A(_03614_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _14598_ (.A0(\fifo0.fifo_store[119][14] ),
    .A1(_06302_),
    .S(_03599_),
    .X(_03615_));
 sky130_fd_sc_hd__clkbuf_1 _14599_ (.A(_03615_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _14600_ (.A0(\fifo0.fifo_store[119][15] ),
    .A1(_06304_),
    .S(_03599_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_1 _14601_ (.A(_03616_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_4 _14602_ (.A(_03964_),
    .B(_04145_),
    .Y(_03617_));
 sky130_fd_sc_hd__buf_8 _14603_ (.A(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _14604_ (.A0(\fifo0.fifo_store[69][0] ),
    .A1(_06283_),
    .S(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _14605_ (.A(_03619_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _14606_ (.A0(\fifo0.fifo_store[69][1] ),
    .A1(_06287_),
    .S(_03618_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _14607_ (.A(_03620_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _14608_ (.A0(\fifo0.fifo_store[69][2] ),
    .A1(_06310_),
    .S(_03618_),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _14609_ (.A(_03621_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _14610_ (.A0(\fifo0.fifo_store[69][3] ),
    .A1(_06312_),
    .S(_03618_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _14611_ (.A(_03622_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _14612_ (.A0(\fifo0.fifo_store[69][4] ),
    .A1(_06314_),
    .S(_03618_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _14613_ (.A(_03623_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _14614_ (.A0(\fifo0.fifo_store[69][5] ),
    .A1(_03884_),
    .S(_03618_),
    .X(_03624_));
 sky130_fd_sc_hd__clkbuf_1 _14615_ (.A(_03624_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _14616_ (.A0(\fifo0.fifo_store[69][6] ),
    .A1(_06317_),
    .S(_03618_),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _14617_ (.A(_03625_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _14618_ (.A0(\fifo0.fifo_store[69][7] ),
    .A1(_03890_),
    .S(_03618_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _14619_ (.A(_03626_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _14620_ (.A0(\fifo0.fifo_store[69][8] ),
    .A1(_06320_),
    .S(_03618_),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _14621_ (.A(_03627_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _14622_ (.A0(\fifo0.fifo_store[69][9] ),
    .A1(_06322_),
    .S(_03618_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _14623_ (.A(_03628_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _14624_ (.A0(\fifo0.fifo_store[69][10] ),
    .A1(_03899_),
    .S(_03617_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _14625_ (.A(_03629_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(\fifo0.fifo_store[69][11] ),
    .A1(_03902_),
    .S(_03617_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _14627_ (.A(_03630_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _14628_ (.A0(\fifo0.fifo_store[69][12] ),
    .A1(_06278_),
    .S(_03617_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _14629_ (.A(_03631_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _14630_ (.A0(\fifo0.fifo_store[69][13] ),
    .A1(_06300_),
    .S(_03617_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _14631_ (.A(_03632_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _14632_ (.A0(\fifo0.fifo_store[69][14] ),
    .A1(_06302_),
    .S(_03617_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _14633_ (.A(_03633_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _14634_ (.A0(\fifo0.fifo_store[69][15] ),
    .A1(_06304_),
    .S(_03617_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_1 _14635_ (.A(_03634_),
    .X(_02068_));
 sky130_fd_sc_hd__inv_2 _14636_ (.A(_03576_),
    .Y(_03635_));
 sky130_fd_sc_hd__a211o_1 _14637_ (.A1(_03564_),
    .A2(_03566_),
    .B1(_03577_),
    .C1(_03562_),
    .X(_03636_));
 sky130_fd_sc_hd__a21o_1 _14638_ (.A1(\dsmod0.accu1[14] ),
    .A2(_03312_),
    .B1(_03573_),
    .X(_03637_));
 sky130_fd_sc_hd__and2_1 _14639_ (.A(\dsmod0.accu1[15] ),
    .B(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__nor2_1 _14640_ (.A(\dsmod0.accu1[15] ),
    .B(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__or2_1 _14641_ (.A(_03638_),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__inv_2 _14642_ (.A(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__a21oi_1 _14643_ (.A1(_03635_),
    .A2(_03636_),
    .B1(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__a31o_1 _14644_ (.A1(_03635_),
    .A2(_03641_),
    .A3(_03636_),
    .B1(_03333_),
    .X(_03643_));
 sky130_fd_sc_hd__o2bb2a_1 _14645_ (.A1_N(\dsmod0.mod2_out[0] ),
    .A2_N(_03334_),
    .B1(_03642_),
    .B2(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__nor2_1 _14646_ (.A(_05924_),
    .B(_03644_),
    .Y(_02069_));
 sky130_fd_sc_hd__o221a_1 _14647_ (.A1(\dsmod0.mod2_out[1] ),
    .A2(_03330_),
    .B1(_03638_),
    .B2(_03643_),
    .C1(_03361_),
    .X(_02070_));
 sky130_fd_sc_hd__nor2_8 _14648_ (.A(_03919_),
    .B(_04629_),
    .Y(_03645_));
 sky130_fd_sc_hd__buf_8 _14649_ (.A(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _14650_ (.A0(\fifo0.fifo_store[47][0] ),
    .A1(_06283_),
    .S(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _14651_ (.A(_03647_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(\fifo0.fifo_store[47][1] ),
    .A1(_06287_),
    .S(_03646_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _14653_ (.A(_03648_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _14654_ (.A0(\fifo0.fifo_store[47][2] ),
    .A1(_06310_),
    .S(_03646_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _14655_ (.A(_03649_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(\fifo0.fifo_store[47][3] ),
    .A1(_06312_),
    .S(_03646_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _14657_ (.A(_03650_),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(\fifo0.fifo_store[47][4] ),
    .A1(_06314_),
    .S(_03646_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _14659_ (.A(_03651_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(\fifo0.fifo_store[47][5] ),
    .A1(_03884_),
    .S(_03646_),
    .X(_03652_));
 sky130_fd_sc_hd__clkbuf_1 _14661_ (.A(_03652_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _14662_ (.A0(\fifo0.fifo_store[47][6] ),
    .A1(_06317_),
    .S(_03646_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_1 _14663_ (.A(_03653_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(\fifo0.fifo_store[47][7] ),
    .A1(_03890_),
    .S(_03646_),
    .X(_03654_));
 sky130_fd_sc_hd__clkbuf_1 _14665_ (.A(_03654_),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(\fifo0.fifo_store[47][8] ),
    .A1(_06320_),
    .S(_03646_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _14667_ (.A(_03655_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _14668_ (.A0(\fifo0.fifo_store[47][9] ),
    .A1(_06322_),
    .S(_03646_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _14669_ (.A(_03656_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_1 _14670_ (.A0(\fifo0.fifo_store[47][10] ),
    .A1(_03899_),
    .S(_03645_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _14671_ (.A(_03657_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _14672_ (.A0(\fifo0.fifo_store[47][11] ),
    .A1(_03902_),
    .S(_03645_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_1 _14673_ (.A(_03658_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _14674_ (.A0(\fifo0.fifo_store[47][12] ),
    .A1(_06278_),
    .S(_03645_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_1 _14675_ (.A(_03659_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _14676_ (.A0(\fifo0.fifo_store[47][13] ),
    .A1(_06300_),
    .S(_03645_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_1 _14677_ (.A(_03660_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _14678_ (.A0(\fifo0.fifo_store[47][14] ),
    .A1(_06302_),
    .S(_03645_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _14679_ (.A(_03661_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _14680_ (.A0(\fifo0.fifo_store[47][15] ),
    .A1(_06304_),
    .S(_03645_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _14681_ (.A(_03662_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_8 _14682_ (.A(_03964_),
    .B(_05788_),
    .Y(_03663_));
 sky130_fd_sc_hd__buf_8 _14683_ (.A(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _14684_ (.A0(\fifo0.fifo_store[29][0] ),
    .A1(_06283_),
    .S(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _14685_ (.A(_03665_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _14686_ (.A0(\fifo0.fifo_store[29][1] ),
    .A1(_06287_),
    .S(_03664_),
    .X(_03666_));
 sky130_fd_sc_hd__clkbuf_1 _14687_ (.A(_03666_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _14688_ (.A0(\fifo0.fifo_store[29][2] ),
    .A1(_06310_),
    .S(_03664_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_1 _14689_ (.A(_03667_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _14690_ (.A0(\fifo0.fifo_store[29][3] ),
    .A1(_06312_),
    .S(_03664_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _14691_ (.A(_03668_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _14692_ (.A0(\fifo0.fifo_store[29][4] ),
    .A1(_06314_),
    .S(_03664_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _14693_ (.A(_03669_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _14694_ (.A0(\fifo0.fifo_store[29][5] ),
    .A1(_03884_),
    .S(_03664_),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _14695_ (.A(_03670_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _14696_ (.A0(\fifo0.fifo_store[29][6] ),
    .A1(_06317_),
    .S(_03664_),
    .X(_03671_));
 sky130_fd_sc_hd__clkbuf_1 _14697_ (.A(_03671_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _14698_ (.A0(\fifo0.fifo_store[29][7] ),
    .A1(_03890_),
    .S(_03664_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _14699_ (.A(_03672_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _14700_ (.A0(\fifo0.fifo_store[29][8] ),
    .A1(_06320_),
    .S(_03664_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _14701_ (.A(_03673_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _14702_ (.A0(\fifo0.fifo_store[29][9] ),
    .A1(_06322_),
    .S(_03664_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_1 _14703_ (.A(_03674_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _14704_ (.A0(\fifo0.fifo_store[29][10] ),
    .A1(_03899_),
    .S(_03663_),
    .X(_03675_));
 sky130_fd_sc_hd__clkbuf_1 _14705_ (.A(_03675_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _14706_ (.A0(\fifo0.fifo_store[29][11] ),
    .A1(_03902_),
    .S(_03663_),
    .X(_03676_));
 sky130_fd_sc_hd__clkbuf_1 _14707_ (.A(_03676_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _14708_ (.A0(\fifo0.fifo_store[29][12] ),
    .A1(_06278_),
    .S(_03663_),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_1 _14709_ (.A(_03677_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _14710_ (.A0(\fifo0.fifo_store[29][13] ),
    .A1(_06300_),
    .S(_03663_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _14711_ (.A(_03678_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _14712_ (.A0(\fifo0.fifo_store[29][14] ),
    .A1(_06302_),
    .S(_03663_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _14713_ (.A(_03679_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _14714_ (.A0(\fifo0.fifo_store[29][15] ),
    .A1(_06304_),
    .S(_03663_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _14715_ (.A(_03680_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_8 _14716_ (.A(_03964_),
    .B(_04297_),
    .Y(_03681_));
 sky130_fd_sc_hd__buf_6 _14717_ (.A(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _14718_ (.A0(\fifo0.fifo_store[109][0] ),
    .A1(_06283_),
    .S(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _14719_ (.A(_03683_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _14720_ (.A0(\fifo0.fifo_store[109][1] ),
    .A1(_06287_),
    .S(_03682_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _14721_ (.A(_03684_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _14722_ (.A0(\fifo0.fifo_store[109][2] ),
    .A1(_06310_),
    .S(_03682_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _14723_ (.A(_03685_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _14724_ (.A0(\fifo0.fifo_store[109][3] ),
    .A1(_06312_),
    .S(_03682_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _14725_ (.A(_03686_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _14726_ (.A0(\fifo0.fifo_store[109][4] ),
    .A1(_06314_),
    .S(_03682_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _14727_ (.A(_03687_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _14728_ (.A0(\fifo0.fifo_store[109][5] ),
    .A1(_03884_),
    .S(_03682_),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _14729_ (.A(_03688_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(\fifo0.fifo_store[109][6] ),
    .A1(_06317_),
    .S(_03682_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _14731_ (.A(_03689_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _14732_ (.A0(\fifo0.fifo_store[109][7] ),
    .A1(_03890_),
    .S(_03682_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _14733_ (.A(_03690_),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _14734_ (.A0(\fifo0.fifo_store[109][8] ),
    .A1(_06320_),
    .S(_03682_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_1 _14735_ (.A(_03691_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _14736_ (.A0(\fifo0.fifo_store[109][9] ),
    .A1(_06322_),
    .S(_03682_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_1 _14737_ (.A(_03692_),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _14738_ (.A0(\fifo0.fifo_store[109][10] ),
    .A1(_03899_),
    .S(_03681_),
    .X(_03693_));
 sky130_fd_sc_hd__clkbuf_1 _14739_ (.A(_03693_),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _14740_ (.A0(\fifo0.fifo_store[109][11] ),
    .A1(_03902_),
    .S(_03681_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_1 _14741_ (.A(_03694_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _14742_ (.A0(\fifo0.fifo_store[109][12] ),
    .A1(_06278_),
    .S(_03681_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _14743_ (.A(_03695_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _14744_ (.A0(\fifo0.fifo_store[109][13] ),
    .A1(_06300_),
    .S(_03681_),
    .X(_03696_));
 sky130_fd_sc_hd__clkbuf_1 _14745_ (.A(_03696_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _14746_ (.A0(\fifo0.fifo_store[109][14] ),
    .A1(_06302_),
    .S(_03681_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_1 _14747_ (.A(_03697_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _14748_ (.A0(\fifo0.fifo_store[109][15] ),
    .A1(_06304_),
    .S(_03681_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _14749_ (.A(_03698_),
    .X(_02118_));
 sky130_fd_sc_hd__nor2_1 _14750_ (.A(_06611_),
    .B(_05936_),
    .Y(_03699_));
 sky130_fd_sc_hd__clkbuf_4 _14751_ (.A(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__a21oi_1 _14752_ (.A1(net24),
    .A2(_03700_),
    .B1(_06399_),
    .Y(_03701_));
 sky130_fd_sc_hd__a311oi_1 _14753_ (.A1(_06399_),
    .A2(net24),
    .A3(_03700_),
    .B1(_03701_),
    .C1(_05924_),
    .Y(_02119_));
 sky130_fd_sc_hd__xor2_1 _14754_ (.A(_06380_),
    .B(net25),
    .X(_03702_));
 sky130_fd_sc_hd__and3_1 _14755_ (.A(_06399_),
    .B(net24),
    .C(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__a21oi_1 _14756_ (.A1(_06399_),
    .A2(net24),
    .B1(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__o21ai_1 _14757_ (.A1(_03703_),
    .A2(_03704_),
    .B1(_03700_),
    .Y(_03705_));
 sky130_fd_sc_hd__o211a_1 _14758_ (.A1(_06380_),
    .A2(_03700_),
    .B1(_03705_),
    .C1(_03361_),
    .X(_02120_));
 sky130_fd_sc_hd__a21oi_1 _14759_ (.A1(_06380_),
    .A2(net25),
    .B1(_03703_),
    .Y(_03706_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(_06398_),
    .B(net26),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _14761_ (.A(_06398_),
    .B(net26),
    .Y(_03708_));
 sky130_fd_sc_hd__or2b_1 _14762_ (.A(_03707_),
    .B_N(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__xnor2_1 _14763_ (.A(_03706_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand2_1 _14764_ (.A(_03700_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__o211a_1 _14765_ (.A1(_06398_),
    .A2(_03700_),
    .B1(_03711_),
    .C1(_03361_),
    .X(_02121_));
 sky130_fd_sc_hd__or2_1 _14766_ (.A(_06378_),
    .B(net27),
    .X(_03712_));
 sky130_fd_sc_hd__nand2_1 _14767_ (.A(_06378_),
    .B(net27),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_1 _14768_ (.A(_03712_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__o21ai_1 _14769_ (.A1(_03706_),
    .A2(_03707_),
    .B1(_03708_),
    .Y(_03715_));
 sky130_fd_sc_hd__xor2_1 _14770_ (.A(_03714_),
    .B(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__nand2_1 _14771_ (.A(_03700_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__o211a_1 _14772_ (.A1(_06378_),
    .A2(_03700_),
    .B1(_03717_),
    .C1(_03361_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_1 _14773_ (.A(_06359_),
    .B(net28),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _14774_ (.A(_06359_),
    .B(net28),
    .Y(_03719_));
 sky130_fd_sc_hd__or2b_1 _14775_ (.A(_03718_),
    .B_N(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__a21boi_2 _14776_ (.A1(_03712_),
    .A2(_03715_),
    .B1_N(_03713_),
    .Y(_03721_));
 sky130_fd_sc_hd__xnor2_1 _14777_ (.A(_03720_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_03700_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__o211a_1 _14779_ (.A1(_06359_),
    .A2(_03700_),
    .B1(_03723_),
    .C1(_03361_),
    .X(_02123_));
 sky130_fd_sc_hd__nand2_1 _14780_ (.A(_06918_),
    .B(_05935_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_1 _14781_ (.A(_06405_),
    .B(net29),
    .Y(_03725_));
 sky130_fd_sc_hd__or2_1 _14782_ (.A(_06405_),
    .B(net29),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_1 _14783_ (.A(_03725_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__o21ai_2 _14784_ (.A1(_03718_),
    .A2(_03721_),
    .B1(_03719_),
    .Y(_03728_));
 sky130_fd_sc_hd__xnor2_1 _14785_ (.A(_03727_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _14786_ (.A(_06370_),
    .B(_03724_),
    .Y(_03730_));
 sky130_fd_sc_hd__o211a_1 _14787_ (.A1(_03724_),
    .A2(_03729_),
    .B1(_03730_),
    .C1(_03361_),
    .X(_02124_));
 sky130_fd_sc_hd__a21o_1 _14788_ (.A1(_06405_),
    .A2(net29),
    .B1(_03728_),
    .X(_03731_));
 sky130_fd_sc_hd__a41o_1 _14789_ (.A1(_06919_),
    .A2(_03699_),
    .A3(_03726_),
    .A4(_03731_),
    .B1(_03799_),
    .X(_03732_));
 sky130_fd_sc_hd__a31o_1 _14790_ (.A1(_03699_),
    .A2(_03726_),
    .A3(_03731_),
    .B1(_06919_),
    .X(_03733_));
 sky130_fd_sc_hd__and2b_1 _14791_ (.A_N(_03732_),
    .B(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _14792_ (.A(_03734_),
    .X(_02125_));
 sky130_fd_sc_hd__nor2_8 _14793_ (.A(_03989_),
    .B(_04690_),
    .Y(_03735_));
 sky130_fd_sc_hd__buf_8 _14794_ (.A(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _14795_ (.A0(\fifo0.fifo_store[50][0] ),
    .A1(_06283_),
    .S(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__clkbuf_1 _14796_ (.A(_03737_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _14797_ (.A0(\fifo0.fifo_store[50][1] ),
    .A1(_06287_),
    .S(_03736_),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _14798_ (.A(_03738_),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _14799_ (.A0(\fifo0.fifo_store[50][2] ),
    .A1(_06310_),
    .S(_03736_),
    .X(_03739_));
 sky130_fd_sc_hd__clkbuf_1 _14800_ (.A(_03739_),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _14801_ (.A0(\fifo0.fifo_store[50][3] ),
    .A1(_06312_),
    .S(_03736_),
    .X(_03740_));
 sky130_fd_sc_hd__clkbuf_1 _14802_ (.A(_03740_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _14803_ (.A0(\fifo0.fifo_store[50][4] ),
    .A1(_06314_),
    .S(_03736_),
    .X(_03741_));
 sky130_fd_sc_hd__clkbuf_1 _14804_ (.A(_03741_),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _14805_ (.A0(\fifo0.fifo_store[50][5] ),
    .A1(_03884_),
    .S(_03736_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _14806_ (.A(_03742_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _14807_ (.A0(\fifo0.fifo_store[50][6] ),
    .A1(_06317_),
    .S(_03736_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_1 _14808_ (.A(_03743_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _14809_ (.A0(\fifo0.fifo_store[50][7] ),
    .A1(_03890_),
    .S(_03736_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _14810_ (.A(_03744_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _14811_ (.A0(\fifo0.fifo_store[50][8] ),
    .A1(_06320_),
    .S(_03736_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _14812_ (.A(_03745_),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _14813_ (.A0(\fifo0.fifo_store[50][9] ),
    .A1(_06322_),
    .S(_03736_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _14814_ (.A(_03746_),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _14815_ (.A0(\fifo0.fifo_store[50][10] ),
    .A1(_03899_),
    .S(_03735_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _14816_ (.A(_03747_),
    .X(_02136_));
 sky130_fd_sc_hd__mux2_1 _14817_ (.A0(\fifo0.fifo_store[50][11] ),
    .A1(_03902_),
    .S(_03735_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _14818_ (.A(_03748_),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _14819_ (.A0(\fifo0.fifo_store[50][12] ),
    .A1(_03905_),
    .S(_03735_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _14820_ (.A(_03749_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _14821_ (.A0(\fifo0.fifo_store[50][13] ),
    .A1(_06300_),
    .S(_03735_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _14822_ (.A(_03750_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(\fifo0.fifo_store[50][14] ),
    .A1(_06302_),
    .S(_03735_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _14824_ (.A(_03751_),
    .X(_02140_));
 sky130_fd_sc_hd__mux2_1 _14825_ (.A0(\fifo0.fifo_store[50][15] ),
    .A1(_06304_),
    .S(_03735_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _14826_ (.A(_03752_),
    .X(_02141_));
 sky130_fd_sc_hd__nor2_8 _14827_ (.A(_04031_),
    .B(_04356_),
    .Y(_03753_));
 sky130_fd_sc_hd__buf_12 _14828_ (.A(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _14829_ (.A0(\fifo0.fifo_store[9][0] ),
    .A1(_03821_),
    .S(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _14830_ (.A(_03755_),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(\fifo0.fifo_store[9][1] ),
    .A1(_03872_),
    .S(_03754_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _14832_ (.A(_03756_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(\fifo0.fifo_store[9][2] ),
    .A1(_06310_),
    .S(_03754_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _14834_ (.A(_03757_),
    .X(_02144_));
 sky130_fd_sc_hd__mux2_1 _14835_ (.A0(\fifo0.fifo_store[9][3] ),
    .A1(_06312_),
    .S(_03754_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _14836_ (.A(_03758_),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _14837_ (.A0(\fifo0.fifo_store[9][4] ),
    .A1(_06314_),
    .S(_03754_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _14838_ (.A(_03759_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(\fifo0.fifo_store[9][5] ),
    .A1(_03884_),
    .S(_03754_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_1 _14840_ (.A(_03760_),
    .X(_02147_));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(\fifo0.fifo_store[9][6] ),
    .A1(_06317_),
    .S(_03754_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _14842_ (.A(_03761_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(\fifo0.fifo_store[9][7] ),
    .A1(_03890_),
    .S(_03754_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _14844_ (.A(_03762_),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(\fifo0.fifo_store[9][8] ),
    .A1(_06320_),
    .S(_03754_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _14846_ (.A(_03763_),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\fifo0.fifo_store[9][9] ),
    .A1(_06322_),
    .S(_03754_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _14848_ (.A(_03764_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(\fifo0.fifo_store[9][10] ),
    .A1(_03899_),
    .S(_03753_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_1 _14850_ (.A(_03765_),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(\fifo0.fifo_store[9][11] ),
    .A1(_03902_),
    .S(_03753_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _14852_ (.A(_03766_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(\fifo0.fifo_store[9][12] ),
    .A1(_03905_),
    .S(_03753_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _14854_ (.A(_03767_),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(\fifo0.fifo_store[9][13] ),
    .A1(_03908_),
    .S(_03753_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _14856_ (.A(_03768_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(\fifo0.fifo_store[9][14] ),
    .A1(_03911_),
    .S(_03753_),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_1 _14858_ (.A(_03769_),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _14859_ (.A0(\fifo0.fifo_store[9][15] ),
    .A1(_03914_),
    .S(_03753_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _14860_ (.A(_03770_),
    .X(_02157_));
 sky130_fd_sc_hd__nor2_1 _14861_ (.A(_05944_),
    .B(_05945_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _14862_ (.A(_05946_),
    .B(_05947_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _14863_ (.A(_05948_),
    .B(_05949_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_1 _14864_ (.A(_05950_),
    .B(_05951_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _14865_ (.A(_05952_),
    .B(_05953_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _14866_ (.A(_05955_),
    .B(_05956_),
    .Y(_02163_));
 sky130_fd_sc_hd__a21oi_1 _14867_ (.A1(\fifo0.read_ptr[6] ),
    .A2(_05955_),
    .B1(_05957_),
    .Y(_02164_));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00007_),
    .Q(\fifo0.fifo_store[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00008_),
    .Q(\fifo0.fifo_store[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00009_),
    .Q(\fifo0.fifo_store[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00010_),
    .Q(\fifo0.fifo_store[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00011_),
    .Q(\fifo0.fifo_store[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_301_clk_i),
    .D(_00012_),
    .Q(\fifo0.fifo_store[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00013_),
    .Q(\fifo0.fifo_store[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00014_),
    .Q(\fifo0.fifo_store[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_302_clk_i),
    .D(_00015_),
    .Q(\fifo0.fifo_store[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00016_),
    .Q(\fifo0.fifo_store[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00017_),
    .Q(\fifo0.fifo_store[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00018_),
    .Q(\fifo0.fifo_store[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00019_),
    .Q(\fifo0.fifo_store[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00020_),
    .Q(\fifo0.fifo_store[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00021_),
    .Q(\fifo0.fifo_store[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00022_),
    .Q(\fifo0.fifo_store[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_60_clk_i),
    .D(_00023_),
    .Q(\fifo0.fifo_store[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_60_clk_i),
    .D(_00024_),
    .Q(\fifo0.fifo_store[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_120_clk_i),
    .D(_00025_),
    .Q(\fifo0.fifo_store[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_49_clk_i),
    .D(_00026_),
    .Q(\fifo0.fifo_store[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_48_clk_i),
    .D(_00027_),
    .Q(\fifo0.fifo_store[80][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_125_clk_i),
    .D(_00028_),
    .Q(\fifo0.fifo_store[80][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_120_clk_i),
    .D(_00029_),
    .Q(\fifo0.fifo_store[80][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00030_),
    .Q(\fifo0.fifo_store[80][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00031_),
    .Q(\fifo0.fifo_store[80][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_42_clk_i),
    .D(_00032_),
    .Q(\fifo0.fifo_store[80][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00033_),
    .Q(\fifo0.fifo_store[80][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00034_),
    .Q(\fifo0.fifo_store[80][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00035_),
    .Q(\fifo0.fifo_store[80][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00036_),
    .Q(\fifo0.fifo_store[80][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00037_),
    .Q(\fifo0.fifo_store[80][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00038_),
    .Q(\fifo0.fifo_store[80][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00039_),
    .Q(\fifo0.fifo_store[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00040_),
    .Q(\fifo0.fifo_store[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_304_clk_i),
    .D(_00041_),
    .Q(\fifo0.fifo_store[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00042_),
    .Q(\fifo0.fifo_store[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00043_),
    .Q(\fifo0.fifo_store[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_303_clk_i),
    .D(_00044_),
    .Q(\fifo0.fifo_store[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00045_),
    .Q(\fifo0.fifo_store[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00046_),
    .Q(\fifo0.fifo_store[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_302_clk_i),
    .D(_00047_),
    .Q(\fifo0.fifo_store[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00048_),
    .Q(\fifo0.fifo_store[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00049_),
    .Q(\fifo0.fifo_store[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00050_),
    .Q(\fifo0.fifo_store[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00051_),
    .Q(\fifo0.fifo_store[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00052_),
    .Q(\fifo0.fifo_store[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00053_),
    .Q(\fifo0.fifo_store[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00054_),
    .Q(\fifo0.fifo_store[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00055_),
    .Q(\fifo0.fifo_store[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00056_),
    .Q(\fifo0.fifo_store[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00057_),
    .Q(\fifo0.fifo_store[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00058_),
    .Q(\fifo0.fifo_store[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00059_),
    .Q(\fifo0.fifo_store[78][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_302_clk_i),
    .D(_00060_),
    .Q(\fifo0.fifo_store[78][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00061_),
    .Q(\fifo0.fifo_store[78][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_300_clk_i),
    .D(_00062_),
    .Q(\fifo0.fifo_store[78][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00063_),
    .Q(\fifo0.fifo_store[78][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00064_),
    .Q(\fifo0.fifo_store[78][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00065_),
    .Q(\fifo0.fifo_store[78][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00066_),
    .Q(\fifo0.fifo_store[78][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00067_),
    .Q(\fifo0.fifo_store[78][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00068_),
    .Q(\fifo0.fifo_store[78][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00069_),
    .Q(\fifo0.fifo_store[78][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00070_),
    .Q(\fifo0.fifo_store[78][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00071_),
    .Q(\fifo0.fifo_store[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_57_clk_i),
    .D(_00072_),
    .Q(\fifo0.fifo_store[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00073_),
    .Q(\fifo0.fifo_store[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00074_),
    .Q(\fifo0.fifo_store[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00075_),
    .Q(\fifo0.fifo_store[77][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_302_clk_i),
    .D(_00076_),
    .Q(\fifo0.fifo_store[77][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00077_),
    .Q(\fifo0.fifo_store[77][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00078_),
    .Q(\fifo0.fifo_store[77][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00079_),
    .Q(\fifo0.fifo_store[77][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00080_),
    .Q(\fifo0.fifo_store[77][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00081_),
    .Q(\fifo0.fifo_store[77][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00082_),
    .Q(\fifo0.fifo_store[77][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00083_),
    .Q(\fifo0.fifo_store[77][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00084_),
    .Q(\fifo0.fifo_store[77][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00085_),
    .Q(\fifo0.fifo_store[77][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00086_),
    .Q(\fifo0.fifo_store[77][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_58_clk_i),
    .D(_00087_),
    .Q(\fifo0.fifo_store[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_58_clk_i),
    .D(_00088_),
    .Q(\fifo0.fifo_store[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00089_),
    .Q(\fifo0.fifo_store[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_54_clk_i),
    .D(_00090_),
    .Q(\fifo0.fifo_store[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00091_),
    .Q(\fifo0.fifo_store[98][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_123_clk_i),
    .D(_00092_),
    .Q(\fifo0.fifo_store[98][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00093_),
    .Q(\fifo0.fifo_store[98][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00094_),
    .Q(\fifo0.fifo_store[98][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_124_clk_i),
    .D(_00095_),
    .Q(\fifo0.fifo_store[98][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00096_),
    .Q(\fifo0.fifo_store[98][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00097_),
    .Q(\fifo0.fifo_store[98][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00098_),
    .Q(\fifo0.fifo_store[98][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_241_clk_i),
    .D(_00099_),
    .Q(\fifo0.fifo_store[98][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00100_),
    .Q(\fifo0.fifo_store[98][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00101_),
    .Q(\fifo0.fifo_store[98][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00102_),
    .Q(\fifo0.fifo_store[98][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14964_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00103_),
    .Q(\fifo0.fifo_store[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00104_),
    .Q(\fifo0.fifo_store[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00105_),
    .Q(\fifo0.fifo_store[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00106_),
    .Q(\fifo0.fifo_store[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14968_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00107_),
    .Q(\fifo0.fifo_store[76][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.CLK(clknet_leaf_302_clk_i),
    .D(_00108_),
    .Q(\fifo0.fifo_store[76][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00109_),
    .Q(\fifo0.fifo_store[76][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00110_),
    .Q(\fifo0.fifo_store[76][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00111_),
    .Q(\fifo0.fifo_store[76][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00112_),
    .Q(\fifo0.fifo_store[76][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00113_),
    .Q(\fifo0.fifo_store[76][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00114_),
    .Q(\fifo0.fifo_store[76][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_241_clk_i),
    .D(_00115_),
    .Q(\fifo0.fifo_store[76][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00116_),
    .Q(\fifo0.fifo_store[76][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00117_),
    .Q(\fifo0.fifo_store[76][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00118_),
    .Q(\fifo0.fifo_store[76][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_58_clk_i),
    .D(_00119_),
    .Q(\fifo0.fifo_store[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_58_clk_i),
    .D(_00120_),
    .Q(\fifo0.fifo_store[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00121_),
    .Q(\fifo0.fifo_store[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00122_),
    .Q(\fifo0.fifo_store[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00123_),
    .Q(\fifo0.fifo_store[97][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.CLK(clknet_leaf_123_clk_i),
    .D(_00124_),
    .Q(\fifo0.fifo_store[97][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00125_),
    .Q(\fifo0.fifo_store[97][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00126_),
    .Q(\fifo0.fifo_store[97][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_125_clk_i),
    .D(_00127_),
    .Q(\fifo0.fifo_store[97][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00128_),
    .Q(\fifo0.fifo_store[97][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00129_),
    .Q(\fifo0.fifo_store[97][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00130_),
    .Q(\fifo0.fifo_store[97][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00131_),
    .Q(\fifo0.fifo_store[97][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00132_),
    .Q(\fifo0.fifo_store[97][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00133_),
    .Q(\fifo0.fifo_store[97][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00134_),
    .Q(\fifo0.fifo_store[97][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00135_),
    .Q(\fifo0.fifo_store[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_57_clk_i),
    .D(_00136_),
    .Q(\fifo0.fifo_store[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00137_),
    .Q(\fifo0.fifo_store[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00138_),
    .Q(\fifo0.fifo_store[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00139_),
    .Q(\fifo0.fifo_store[75][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00140_),
    .Q(\fifo0.fifo_store[75][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00141_),
    .Q(\fifo0.fifo_store[75][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00142_),
    .Q(\fifo0.fifo_store[75][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_300_clk_i),
    .D(_00143_),
    .Q(\fifo0.fifo_store[75][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00144_),
    .Q(\fifo0.fifo_store[75][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00145_),
    .Q(\fifo0.fifo_store[75][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00146_),
    .Q(\fifo0.fifo_store[75][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00147_),
    .Q(\fifo0.fifo_store[75][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00148_),
    .Q(\fifo0.fifo_store[75][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00149_),
    .Q(\fifo0.fifo_store[75][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00150_),
    .Q(\fifo0.fifo_store[75][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_57_clk_i),
    .D(_00151_),
    .Q(\fifo0.fifo_store[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_58_clk_i),
    .D(_00152_),
    .Q(\fifo0.fifo_store[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00153_),
    .Q(\fifo0.fifo_store[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_54_clk_i),
    .D(_00154_),
    .Q(\fifo0.fifo_store[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00155_),
    .Q(\fifo0.fifo_store[96][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_124_clk_i),
    .D(_00156_),
    .Q(\fifo0.fifo_store[96][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00157_),
    .Q(\fifo0.fifo_store[96][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00158_),
    .Q(\fifo0.fifo_store[96][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.CLK(clknet_leaf_125_clk_i),
    .D(_00159_),
    .Q(\fifo0.fifo_store[96][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00160_),
    .Q(\fifo0.fifo_store[96][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00161_),
    .Q(\fifo0.fifo_store[96][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00162_),
    .Q(\fifo0.fifo_store[96][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00163_),
    .Q(\fifo0.fifo_store[96][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00164_),
    .Q(\fifo0.fifo_store[96][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00165_),
    .Q(\fifo0.fifo_store[96][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00166_),
    .Q(\fifo0.fifo_store[96][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00167_),
    .Q(\fifo0.fifo_store[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00168_),
    .Q(\fifo0.fifo_store[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00169_),
    .Q(\fifo0.fifo_store[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00170_),
    .Q(\fifo0.fifo_store[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00171_),
    .Q(\fifo0.fifo_store[74][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00172_),
    .Q(\fifo0.fifo_store[74][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00173_),
    .Q(\fifo0.fifo_store[74][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00174_),
    .Q(\fifo0.fifo_store[74][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_301_clk_i),
    .D(_00175_),
    .Q(\fifo0.fifo_store[74][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00176_),
    .Q(\fifo0.fifo_store[74][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00177_),
    .Q(\fifo0.fifo_store[74][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00178_),
    .Q(\fifo0.fifo_store[74][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00179_),
    .Q(\fifo0.fifo_store[74][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15041_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00180_),
    .Q(\fifo0.fifo_store[74][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00181_),
    .Q(\fifo0.fifo_store[74][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00182_),
    .Q(\fifo0.fifo_store[74][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00183_),
    .Q(\fifo0.fifo_store[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15045_ (.CLK(clknet_leaf_57_clk_i),
    .D(_00184_),
    .Q(\fifo0.fifo_store[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00185_),
    .Q(\fifo0.fifo_store[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00186_),
    .Q(\fifo0.fifo_store[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.CLK(clknet_leaf_53_clk_i),
    .D(_00187_),
    .Q(\fifo0.fifo_store[73][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00188_),
    .Q(\fifo0.fifo_store[73][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00189_),
    .Q(\fifo0.fifo_store[73][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00190_),
    .Q(\fifo0.fifo_store[73][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.CLK(clknet_leaf_300_clk_i),
    .D(_00191_),
    .Q(\fifo0.fifo_store[73][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00192_),
    .Q(\fifo0.fifo_store[73][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00193_),
    .Q(\fifo0.fifo_store[73][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00194_),
    .Q(\fifo0.fifo_store[73][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00195_),
    .Q(\fifo0.fifo_store[73][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00196_),
    .Q(\fifo0.fifo_store[73][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00197_),
    .Q(\fifo0.fifo_store[73][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00198_),
    .Q(\fifo0.fifo_store[73][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00199_),
    .Q(\fifo0.fifo_store[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.CLK(clknet_leaf_57_clk_i),
    .D(_00200_),
    .Q(\fifo0.fifo_store[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.CLK(clknet_leaf_321_clk_i),
    .D(_00201_),
    .Q(\fifo0.fifo_store[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00202_),
    .Q(\fifo0.fifo_store[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00203_),
    .Q(\fifo0.fifo_store[72][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00204_),
    .Q(\fifo0.fifo_store[72][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.CLK(clknet_leaf_320_clk_i),
    .D(_00205_),
    .Q(\fifo0.fifo_store[72][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15067_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00206_),
    .Q(\fifo0.fifo_store[72][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.CLK(clknet_leaf_301_clk_i),
    .D(_00207_),
    .Q(\fifo0.fifo_store[72][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00208_),
    .Q(\fifo0.fifo_store[72][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00209_),
    .Q(\fifo0.fifo_store[72][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00210_),
    .Q(\fifo0.fifo_store[72][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00211_),
    .Q(\fifo0.fifo_store[72][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00212_),
    .Q(\fifo0.fifo_store[72][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15074_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00213_),
    .Q(\fifo0.fifo_store[72][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00214_),
    .Q(\fifo0.fifo_store[72][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_62_clk_i),
    .D(_00215_),
    .Q(\fifo0.fifo_store[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.CLK(clknet_leaf_59_clk_i),
    .D(_00216_),
    .Q(\fifo0.fifo_store[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00217_),
    .Q(\fifo0.fifo_store[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.CLK(clknet_leaf_61_clk_i),
    .D(_00218_),
    .Q(\fifo0.fifo_store[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.CLK(clknet_leaf_50_clk_i),
    .D(_00219_),
    .Q(\fifo0.fifo_store[71][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00220_),
    .Q(\fifo0.fifo_store[71][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.CLK(clknet_leaf_116_clk_i),
    .D(_00221_),
    .Q(\fifo0.fifo_store[71][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00222_),
    .Q(\fifo0.fifo_store[71][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.CLK(clknet_leaf_127_clk_i),
    .D(_00223_),
    .Q(\fifo0.fifo_store[71][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00224_),
    .Q(\fifo0.fifo_store[71][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00225_),
    .Q(\fifo0.fifo_store[71][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00226_),
    .Q(\fifo0.fifo_store[71][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00227_),
    .Q(\fifo0.fifo_store[71][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00228_),
    .Q(\fifo0.fifo_store[71][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00229_),
    .Q(\fifo0.fifo_store[71][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00230_),
    .Q(\fifo0.fifo_store[71][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00231_),
    .Q(\fifo0.fifo_store[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_81_clk_i),
    .D(_00232_),
    .Q(\fifo0.fifo_store[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_112_clk_i),
    .D(_00233_),
    .Q(\fifo0.fifo_store[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.CLK(clknet_leaf_70_clk_i),
    .D(_00234_),
    .Q(\fifo0.fifo_store[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00235_),
    .Q(\fifo0.fifo_store[95][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00236_),
    .Q(\fifo0.fifo_store[95][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.CLK(clknet_leaf_117_clk_i),
    .D(_00237_),
    .Q(\fifo0.fifo_store[95][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00238_),
    .Q(\fifo0.fifo_store[95][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.CLK(clknet_leaf_135_clk_i),
    .D(_00239_),
    .Q(\fifo0.fifo_store[95][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.CLK(clknet_leaf_113_clk_i),
    .D(_00240_),
    .Q(\fifo0.fifo_store[95][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00241_),
    .Q(\fifo0.fifo_store[95][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00242_),
    .Q(\fifo0.fifo_store[95][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00243_),
    .Q(\fifo0.fifo_store[95][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00244_),
    .Q(\fifo0.fifo_store[95][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00245_),
    .Q(\fifo0.fifo_store[95][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_159_clk_i),
    .D(_00246_),
    .Q(\fifo0.fifo_store[95][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_62_clk_i),
    .D(_00247_),
    .Q(\fifo0.fifo_store[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_59_clk_i),
    .D(_00248_),
    .Q(\fifo0.fifo_store[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_121_clk_i),
    .D(_00249_),
    .Q(\fifo0.fifo_store[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_62_clk_i),
    .D(_00250_),
    .Q(\fifo0.fifo_store[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_50_clk_i),
    .D(_00251_),
    .Q(\fifo0.fifo_store[70][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00252_),
    .Q(\fifo0.fifo_store[70][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_115_clk_i),
    .D(_00253_),
    .Q(\fifo0.fifo_store[70][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00254_),
    .Q(\fifo0.fifo_store[70][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_126_clk_i),
    .D(_00255_),
    .Q(\fifo0.fifo_store[70][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_42_clk_i),
    .D(_00256_),
    .Q(\fifo0.fifo_store[70][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00257_),
    .Q(\fifo0.fifo_store[70][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00258_),
    .Q(\fifo0.fifo_store[70][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00259_),
    .Q(\fifo0.fifo_store[70][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00260_),
    .Q(\fifo0.fifo_store[70][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00261_),
    .Q(\fifo0.fifo_store[70][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00262_),
    .Q(\fifo0.fifo_store[70][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15124_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00263_),
    .Q(\fifo0.fifo_store[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00264_),
    .Q(\fifo0.fifo_store[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00265_),
    .Q(\fifo0.fifo_store[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00266_),
    .Q(\fifo0.fifo_store[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00267_),
    .Q(\fifo0.fifo_store[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.CLK(clknet_leaf_303_clk_i),
    .D(_00268_),
    .Q(\fifo0.fifo_store[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00269_),
    .Q(\fifo0.fifo_store[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00270_),
    .Q(\fifo0.fifo_store[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00271_),
    .Q(\fifo0.fifo_store[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00272_),
    .Q(\fifo0.fifo_store[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00273_),
    .Q(\fifo0.fifo_store[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15135_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00274_),
    .Q(\fifo0.fifo_store[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15136_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00275_),
    .Q(\fifo0.fifo_store[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15137_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00276_),
    .Q(\fifo0.fifo_store[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15138_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00277_),
    .Q(\fifo0.fifo_store[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15139_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00278_),
    .Q(\fifo0.fifo_store[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15140_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00279_),
    .Q(\fifo0.fifo_store[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.CLK(clknet_leaf_81_clk_i),
    .D(_00280_),
    .Q(\fifo0.fifo_store[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.CLK(clknet_leaf_109_clk_i),
    .D(_00281_),
    .Q(\fifo0.fifo_store[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00282_),
    .Q(\fifo0.fifo_store[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00283_),
    .Q(\fifo0.fifo_store[93][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00284_),
    .Q(\fifo0.fifo_store[93][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00285_),
    .Q(\fifo0.fifo_store[93][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00286_),
    .Q(\fifo0.fifo_store[93][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.CLK(clknet_leaf_135_clk_i),
    .D(_00287_),
    .Q(\fifo0.fifo_store[93][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.CLK(clknet_leaf_113_clk_i),
    .D(_00288_),
    .Q(\fifo0.fifo_store[93][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.CLK(clknet_leaf_159_clk_i),
    .D(_00289_),
    .Q(\fifo0.fifo_store[93][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00290_),
    .Q(\fifo0.fifo_store[93][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00291_),
    .Q(\fifo0.fifo_store[93][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15153_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00292_),
    .Q(\fifo0.fifo_store[93][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15154_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00293_),
    .Q(\fifo0.fifo_store[93][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15155_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00294_),
    .Q(\fifo0.fifo_store[93][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15156_ (.CLK(clknet_leaf_62_clk_i),
    .D(_00295_),
    .Q(\fifo0.fifo_store[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15157_ (.CLK(clknet_leaf_59_clk_i),
    .D(_00296_),
    .Q(\fifo0.fifo_store[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15158_ (.CLK(clknet_leaf_121_clk_i),
    .D(_00297_),
    .Q(\fifo0.fifo_store[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15159_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00298_),
    .Q(\fifo0.fifo_store[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15160_ (.CLK(clknet_leaf_51_clk_i),
    .D(_00299_),
    .Q(\fifo0.fifo_store[68][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15161_ (.CLK(clknet_leaf_129_clk_i),
    .D(_00300_),
    .Q(\fifo0.fifo_store[68][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15162_ (.CLK(clknet_leaf_116_clk_i),
    .D(_00301_),
    .Q(\fifo0.fifo_store[68][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15163_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00302_),
    .Q(\fifo0.fifo_store[68][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15164_ (.CLK(clknet_leaf_126_clk_i),
    .D(_00303_),
    .Q(\fifo0.fifo_store[68][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15165_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00304_),
    .Q(\fifo0.fifo_store[68][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15166_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00305_),
    .Q(\fifo0.fifo_store[68][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15167_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00306_),
    .Q(\fifo0.fifo_store[68][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15168_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00307_),
    .Q(\fifo0.fifo_store[68][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15169_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00308_),
    .Q(\fifo0.fifo_store[68][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15170_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00309_),
    .Q(\fifo0.fifo_store[68][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15171_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00310_),
    .Q(\fifo0.fifo_store[68][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15172_ (.CLK(clknet_leaf_69_clk_i),
    .D(_00311_),
    .Q(\fifo0.fifo_store[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15173_ (.CLK(clknet_leaf_81_clk_i),
    .D(_00312_),
    .Q(\fifo0.fifo_store[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15174_ (.CLK(clknet_leaf_109_clk_i),
    .D(_00313_),
    .Q(\fifo0.fifo_store[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15175_ (.CLK(clknet_leaf_70_clk_i),
    .D(_00314_),
    .Q(\fifo0.fifo_store[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15176_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00315_),
    .Q(\fifo0.fifo_store[92][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15177_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00316_),
    .Q(\fifo0.fifo_store[92][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15178_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00317_),
    .Q(\fifo0.fifo_store[92][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15179_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00318_),
    .Q(\fifo0.fifo_store[92][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15180_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00319_),
    .Q(\fifo0.fifo_store[92][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15181_ (.CLK(clknet_leaf_113_clk_i),
    .D(_00320_),
    .Q(\fifo0.fifo_store[92][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15182_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00321_),
    .Q(\fifo0.fifo_store[92][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15183_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00322_),
    .Q(\fifo0.fifo_store[92][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15184_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00323_),
    .Q(\fifo0.fifo_store[92][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15185_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00324_),
    .Q(\fifo0.fifo_store[92][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15186_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00325_),
    .Q(\fifo0.fifo_store[92][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15187_ (.CLK(clknet_leaf_159_clk_i),
    .D(_00326_),
    .Q(\fifo0.fifo_store[92][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15188_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00327_),
    .Q(\fifo0.fifo_store[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15189_ (.CLK(clknet_leaf_79_clk_i),
    .D(_00328_),
    .Q(\fifo0.fifo_store[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15190_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00329_),
    .Q(\fifo0.fifo_store[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15191_ (.CLK(clknet_leaf_68_clk_i),
    .D(_00330_),
    .Q(\fifo0.fifo_store[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15192_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00331_),
    .Q(\fifo0.fifo_store[105][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15193_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00332_),
    .Q(\fifo0.fifo_store[105][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15194_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00333_),
    .Q(\fifo0.fifo_store[105][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15195_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00334_),
    .Q(\fifo0.fifo_store[105][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15196_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00335_),
    .Q(\fifo0.fifo_store[105][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15197_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00336_),
    .Q(\fifo0.fifo_store[105][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15198_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00337_),
    .Q(\fifo0.fifo_store[105][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15199_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00338_),
    .Q(\fifo0.fifo_store[105][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15200_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00339_),
    .Q(\fifo0.fifo_store[105][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15201_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00340_),
    .Q(\fifo0.fifo_store[105][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15202_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00341_),
    .Q(\fifo0.fifo_store[105][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00342_),
    .Q(\fifo0.fifo_store[105][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00343_),
    .Q(\fifo0.fifo_store[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15205_ (.CLK(clknet_leaf_72_clk_i),
    .D(_00344_),
    .Q(\fifo0.fifo_store[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.CLK(clknet_leaf_110_clk_i),
    .D(_00345_),
    .Q(\fifo0.fifo_store[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15207_ (.CLK(clknet_leaf_72_clk_i),
    .D(_00346_),
    .Q(\fifo0.fifo_store[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00347_),
    .Q(\fifo0.fifo_store[118][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15209_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00348_),
    .Q(\fifo0.fifo_store[118][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15210_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00349_),
    .Q(\fifo0.fifo_store[118][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15211_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00350_),
    .Q(\fifo0.fifo_store[118][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15212_ (.CLK(clknet_leaf_141_clk_i),
    .D(_00351_),
    .Q(\fifo0.fifo_store[118][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15213_ (.CLK(clknet_leaf_112_clk_i),
    .D(_00352_),
    .Q(\fifo0.fifo_store[118][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15214_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00353_),
    .Q(\fifo0.fifo_store[118][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15215_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00354_),
    .Q(\fifo0.fifo_store[118][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00355_),
    .Q(\fifo0.fifo_store[118][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00356_),
    .Q(\fifo0.fifo_store[118][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15218_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00357_),
    .Q(\fifo0.fifo_store[118][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15219_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00358_),
    .Q(\fifo0.fifo_store[118][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15220_ (.CLK(clknet_leaf_78_clk_i),
    .D(_00359_),
    .Q(\fifo0.fifo_store[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15221_ (.CLK(clknet_leaf_78_clk_i),
    .D(_00360_),
    .Q(\fifo0.fifo_store[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15222_ (.CLK(clknet_leaf_104_clk_i),
    .D(_00361_),
    .Q(\fifo0.fifo_store[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15223_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00362_),
    .Q(\fifo0.fifo_store[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15224_ (.CLK(clknet_leaf_84_clk_i),
    .D(_00363_),
    .Q(\fifo0.fifo_store[115][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15225_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00364_),
    .Q(\fifo0.fifo_store[115][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15226_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00365_),
    .Q(\fifo0.fifo_store[115][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15227_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00366_),
    .Q(\fifo0.fifo_store[115][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15228_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00367_),
    .Q(\fifo0.fifo_store[115][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00368_),
    .Q(\fifo0.fifo_store[115][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00369_),
    .Q(\fifo0.fifo_store[115][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00370_),
    .Q(\fifo0.fifo_store[115][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00371_),
    .Q(\fifo0.fifo_store[115][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00372_),
    .Q(\fifo0.fifo_store[115][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00373_),
    .Q(\fifo0.fifo_store[115][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00374_),
    .Q(\fifo0.fifo_store[115][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.CLK(clknet_leaf_61_clk_i),
    .D(_00375_),
    .Q(\fifo0.fifo_store[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.CLK(clknet_leaf_81_clk_i),
    .D(_00376_),
    .Q(\fifo0.fifo_store[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15238_ (.CLK(clknet_leaf_91_clk_i),
    .D(_00377_),
    .Q(\fifo0.fifo_store[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00378_),
    .Q(\fifo0.fifo_store[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.CLK(clknet_leaf_84_clk_i),
    .D(_00379_),
    .Q(\fifo0.fifo_store[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00380_),
    .Q(\fifo0.fifo_store[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00381_),
    .Q(\fifo0.fifo_store[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00382_),
    .Q(\fifo0.fifo_store[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00383_),
    .Q(\fifo0.fifo_store[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00384_),
    .Q(\fifo0.fifo_store[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00385_),
    .Q(\fifo0.fifo_store[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00386_),
    .Q(\fifo0.fifo_store[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00387_),
    .Q(\fifo0.fifo_store[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00388_),
    .Q(\fifo0.fifo_store[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00389_),
    .Q(\fifo0.fifo_store[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15251_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00390_),
    .Q(\fifo0.fifo_store[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15252_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00391_),
    .Q(\fifo0.fifo_store[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15253_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00392_),
    .Q(\fifo0.fifo_store[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15254_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00393_),
    .Q(\fifo0.fifo_store[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15255_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00394_),
    .Q(\fifo0.fifo_store[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00395_),
    .Q(\fifo0.fifo_store[120][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00396_),
    .Q(\fifo0.fifo_store[120][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00397_),
    .Q(\fifo0.fifo_store[120][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00398_),
    .Q(\fifo0.fifo_store[120][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00399_),
    .Q(\fifo0.fifo_store[120][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00400_),
    .Q(\fifo0.fifo_store[120][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00401_),
    .Q(\fifo0.fifo_store[120][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00402_),
    .Q(\fifo0.fifo_store[120][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00403_),
    .Q(\fifo0.fifo_store[120][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00404_),
    .Q(\fifo0.fifo_store[120][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00405_),
    .Q(\fifo0.fifo_store[120][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00406_),
    .Q(\fifo0.fifo_store[120][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00407_),
    .Q(\fifo0.fifo_store[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15269_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00408_),
    .Q(\fifo0.fifo_store[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15270_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00409_),
    .Q(\fifo0.fifo_store[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00410_),
    .Q(\fifo0.fifo_store[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00411_),
    .Q(\fifo0.fifo_store[121][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00412_),
    .Q(\fifo0.fifo_store[121][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00413_),
    .Q(\fifo0.fifo_store[121][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15275_ (.CLK(clknet_leaf_149_clk_i),
    .D(_00414_),
    .Q(\fifo0.fifo_store[121][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00415_),
    .Q(\fifo0.fifo_store[121][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00416_),
    .Q(\fifo0.fifo_store[121][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00417_),
    .Q(\fifo0.fifo_store[121][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00418_),
    .Q(\fifo0.fifo_store[121][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00419_),
    .Q(\fifo0.fifo_store[121][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00420_),
    .Q(\fifo0.fifo_store[121][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15282_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00421_),
    .Q(\fifo0.fifo_store[121][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00422_),
    .Q(\fifo0.fifo_store[121][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00423_),
    .Q(\fifo0.fifo_store[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00424_),
    .Q(\fifo0.fifo_store[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00425_),
    .Q(\fifo0.fifo_store[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00426_),
    .Q(\fifo0.fifo_store[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00427_),
    .Q(\fifo0.fifo_store[122][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15289_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00428_),
    .Q(\fifo0.fifo_store[122][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00429_),
    .Q(\fifo0.fifo_store[122][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00430_),
    .Q(\fifo0.fifo_store[122][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15292_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00431_),
    .Q(\fifo0.fifo_store[122][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00432_),
    .Q(\fifo0.fifo_store[122][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00433_),
    .Q(\fifo0.fifo_store[122][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00434_),
    .Q(\fifo0.fifo_store[122][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00435_),
    .Q(\fifo0.fifo_store[122][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00436_),
    .Q(\fifo0.fifo_store[122][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00437_),
    .Q(\fifo0.fifo_store[122][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00438_),
    .Q(\fifo0.fifo_store[122][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.CLK(clknet_leaf_70_clk_i),
    .D(_00439_),
    .Q(\fifo0.fifo_store[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.CLK(clknet_leaf_78_clk_i),
    .D(_00440_),
    .Q(\fifo0.fifo_store[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.CLK(clknet_leaf_105_clk_i),
    .D(_00441_),
    .Q(\fifo0.fifo_store[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00442_),
    .Q(\fifo0.fifo_store[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.CLK(clknet_leaf_85_clk_i),
    .D(_00443_),
    .Q(\fifo0.fifo_store[116][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00444_),
    .Q(\fifo0.fifo_store[116][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.CLK(clknet_leaf_91_clk_i),
    .D(_00445_),
    .Q(\fifo0.fifo_store[116][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00446_),
    .Q(\fifo0.fifo_store[116][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00447_),
    .Q(\fifo0.fifo_store[116][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15309_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00448_),
    .Q(\fifo0.fifo_store[116][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15310_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00449_),
    .Q(\fifo0.fifo_store[116][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15311_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00450_),
    .Q(\fifo0.fifo_store[116][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00451_),
    .Q(\fifo0.fifo_store[116][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00452_),
    .Q(\fifo0.fifo_store[116][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15314_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00453_),
    .Q(\fifo0.fifo_store[116][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15315_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00454_),
    .Q(\fifo0.fifo_store[116][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00455_),
    .Q(\fifo0.fifo_store[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00456_),
    .Q(\fifo0.fifo_store[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00457_),
    .Q(\fifo0.fifo_store[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.CLK(clknet_leaf_82_clk_i),
    .D(_00458_),
    .Q(\fifo0.fifo_store[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.CLK(clknet_leaf_83_clk_i),
    .D(_00459_),
    .Q(\fifo0.fifo_store[123][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00460_),
    .Q(\fifo0.fifo_store[123][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15322_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00461_),
    .Q(\fifo0.fifo_store[123][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15323_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00462_),
    .Q(\fifo0.fifo_store[123][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15324_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00463_),
    .Q(\fifo0.fifo_store[123][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00464_),
    .Q(\fifo0.fifo_store[123][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15326_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00465_),
    .Q(\fifo0.fifo_store[123][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15327_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00466_),
    .Q(\fifo0.fifo_store[123][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15328_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00467_),
    .Q(\fifo0.fifo_store[123][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15329_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00468_),
    .Q(\fifo0.fifo_store[123][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15330_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00469_),
    .Q(\fifo0.fifo_store[123][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15331_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00470_),
    .Q(\fifo0.fifo_store[123][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.CLK(clknet_leaf_70_clk_i),
    .D(_00471_),
    .Q(\fifo0.fifo_store[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15333_ (.CLK(clknet_leaf_77_clk_i),
    .D(_00472_),
    .Q(\fifo0.fifo_store[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15334_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00473_),
    .Q(\fifo0.fifo_store[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15335_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00474_),
    .Q(\fifo0.fifo_store[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.CLK(clknet_leaf_85_clk_i),
    .D(_00475_),
    .Q(\fifo0.fifo_store[117][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15337_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00476_),
    .Q(\fifo0.fifo_store[117][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15338_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00477_),
    .Q(\fifo0.fifo_store[117][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15339_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00478_),
    .Q(\fifo0.fifo_store[117][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15340_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00479_),
    .Q(\fifo0.fifo_store[117][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15341_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00480_),
    .Q(\fifo0.fifo_store[117][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15342_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00481_),
    .Q(\fifo0.fifo_store[117][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15343_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00482_),
    .Q(\fifo0.fifo_store[117][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15344_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00483_),
    .Q(\fifo0.fifo_store[117][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15345_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00484_),
    .Q(\fifo0.fifo_store[117][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15346_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00485_),
    .Q(\fifo0.fifo_store[117][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15347_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00486_),
    .Q(\fifo0.fifo_store[117][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15348_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00487_),
    .Q(\fifo0.fifo_store[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15349_ (.CLK(clknet_leaf_70_clk_i),
    .D(_00488_),
    .Q(\fifo0.fifo_store[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15350_ (.CLK(clknet_leaf_109_clk_i),
    .D(_00489_),
    .Q(\fifo0.fifo_store[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15351_ (.CLK(clknet_leaf_68_clk_i),
    .D(_00490_),
    .Q(\fifo0.fifo_store[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00491_),
    .Q(\fifo0.fifo_store[124][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15353_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00492_),
    .Q(\fifo0.fifo_store[124][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.CLK(clknet_leaf_112_clk_i),
    .D(_00493_),
    .Q(\fifo0.fifo_store[124][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00494_),
    .Q(\fifo0.fifo_store[124][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00495_),
    .Q(\fifo0.fifo_store[124][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.CLK(clknet_leaf_89_clk_i),
    .D(_00496_),
    .Q(\fifo0.fifo_store[124][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15358_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00497_),
    .Q(\fifo0.fifo_store[124][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00498_),
    .Q(\fifo0.fifo_store[124][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00499_),
    .Q(\fifo0.fifo_store[124][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15361_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00500_),
    .Q(\fifo0.fifo_store[124][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15362_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00501_),
    .Q(\fifo0.fifo_store[124][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00502_),
    .Q(\fifo0.fifo_store[124][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.CLK(clknet_leaf_75_clk_i),
    .D(_00503_),
    .Q(\fifo0.fifo_store[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00504_),
    .Q(\fifo0.fifo_store[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.CLK(clknet_leaf_103_clk_i),
    .D(_00505_),
    .Q(\fifo0.fifo_store[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15367_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00506_),
    .Q(\fifo0.fifo_store[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00507_),
    .Q(\fifo0.fifo_store[67][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.CLK(clknet_leaf_103_clk_i),
    .D(_00508_),
    .Q(\fifo0.fifo_store[67][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_91_clk_i),
    .D(_00509_),
    .Q(\fifo0.fifo_store[67][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00510_),
    .Q(\fifo0.fifo_store[67][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00511_),
    .Q(\fifo0.fifo_store[67][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00512_),
    .Q(\fifo0.fifo_store[67][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00513_),
    .Q(\fifo0.fifo_store[67][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00514_),
    .Q(\fifo0.fifo_store[67][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00515_),
    .Q(\fifo0.fifo_store[67][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00516_),
    .Q(\fifo0.fifo_store[67][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00517_),
    .Q(\fifo0.fifo_store[67][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15379_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00518_),
    .Q(\fifo0.fifo_store[67][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00519_),
    .Q(\fifo0.fifo_store[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00520_),
    .Q(\fifo0.fifo_store[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.CLK(clknet_leaf_102_clk_i),
    .D(_00521_),
    .Q(\fifo0.fifo_store[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00522_),
    .Q(\fifo0.fifo_store[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.CLK(clknet_leaf_84_clk_i),
    .D(_00523_),
    .Q(\fifo0.fifo_store[112][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00524_),
    .Q(\fifo0.fifo_store[112][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15386_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00525_),
    .Q(\fifo0.fifo_store[112][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15387_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00526_),
    .Q(\fifo0.fifo_store[112][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15388_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00527_),
    .Q(\fifo0.fifo_store[112][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00528_),
    .Q(\fifo0.fifo_store[112][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00529_),
    .Q(\fifo0.fifo_store[112][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15391_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00530_),
    .Q(\fifo0.fifo_store[112][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00531_),
    .Q(\fifo0.fifo_store[112][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00532_),
    .Q(\fifo0.fifo_store[112][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00533_),
    .Q(\fifo0.fifo_store[112][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00534_),
    .Q(\fifo0.fifo_store[112][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00535_),
    .Q(\fifo0.fifo_store[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15397_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00536_),
    .Q(\fifo0.fifo_store[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15398_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00537_),
    .Q(\fifo0.fifo_store[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15399_ (.CLK(clknet_leaf_75_clk_i),
    .D(_00538_),
    .Q(\fifo0.fifo_store[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15400_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00539_),
    .Q(\fifo0.fifo_store[100][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15401_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00540_),
    .Q(\fifo0.fifo_store[100][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.CLK(clknet_leaf_111_clk_i),
    .D(_00541_),
    .Q(\fifo0.fifo_store[100][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00542_),
    .Q(\fifo0.fifo_store[100][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00543_),
    .Q(\fifo0.fifo_store[100][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15405_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00544_),
    .Q(\fifo0.fifo_store[100][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15406_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00545_),
    .Q(\fifo0.fifo_store[100][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15407_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00546_),
    .Q(\fifo0.fifo_store[100][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15408_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00547_),
    .Q(\fifo0.fifo_store[100][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15409_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00548_),
    .Q(\fifo0.fifo_store[100][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15410_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00549_),
    .Q(\fifo0.fifo_store[100][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15411_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00550_),
    .Q(\fifo0.fifo_store[100][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15412_ (.CLK(clknet_leaf_77_clk_i),
    .D(_00551_),
    .Q(\fifo0.fifo_store[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15413_ (.CLK(clknet_leaf_79_clk_i),
    .D(_00552_),
    .Q(\fifo0.fifo_store[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15414_ (.CLK(clknet_leaf_102_clk_i),
    .D(_00553_),
    .Q(\fifo0.fifo_store[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15415_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00554_),
    .Q(\fifo0.fifo_store[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15416_ (.CLK(clknet_leaf_85_clk_i),
    .D(_00555_),
    .Q(\fifo0.fifo_store[113][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15417_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00556_),
    .Q(\fifo0.fifo_store[113][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15418_ (.CLK(clknet_leaf_91_clk_i),
    .D(_00557_),
    .Q(\fifo0.fifo_store[113][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15419_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00558_),
    .Q(\fifo0.fifo_store[113][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15420_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00559_),
    .Q(\fifo0.fifo_store[113][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15421_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00560_),
    .Q(\fifo0.fifo_store[113][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00561_),
    .Q(\fifo0.fifo_store[113][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15423_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00562_),
    .Q(\fifo0.fifo_store[113][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15424_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00563_),
    .Q(\fifo0.fifo_store[113][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15425_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00564_),
    .Q(\fifo0.fifo_store[113][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15426_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00565_),
    .Q(\fifo0.fifo_store[113][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15427_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00566_),
    .Q(\fifo0.fifo_store[113][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15428_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00567_),
    .Q(\fifo0.fifo_store[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15429_ (.CLK(clknet_leaf_73_clk_i),
    .D(_00568_),
    .Q(\fifo0.fifo_store[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15430_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00569_),
    .Q(\fifo0.fifo_store[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15431_ (.CLK(clknet_leaf_68_clk_i),
    .D(_00570_),
    .Q(\fifo0.fifo_store[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15432_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00571_),
    .Q(\fifo0.fifo_store[111][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15433_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00572_),
    .Q(\fifo0.fifo_store[111][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15434_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00573_),
    .Q(\fifo0.fifo_store[111][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15435_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00574_),
    .Q(\fifo0.fifo_store[111][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15436_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00575_),
    .Q(\fifo0.fifo_store[111][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15437_ (.CLK(clknet_leaf_88_clk_i),
    .D(_00576_),
    .Q(\fifo0.fifo_store[111][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15438_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00577_),
    .Q(\fifo0.fifo_store[111][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15439_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00578_),
    .Q(\fifo0.fifo_store[111][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15440_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00579_),
    .Q(\fifo0.fifo_store[111][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15441_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00580_),
    .Q(\fifo0.fifo_store[111][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00581_),
    .Q(\fifo0.fifo_store[111][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15443_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00582_),
    .Q(\fifo0.fifo_store[111][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.CLK(clknet_leaf_77_clk_i),
    .D(_00583_),
    .Q(\fifo0.fifo_store[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15445_ (.CLK(clknet_leaf_79_clk_i),
    .D(_00584_),
    .Q(\fifo0.fifo_store[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15446_ (.CLK(clknet_leaf_104_clk_i),
    .D(_00585_),
    .Q(\fifo0.fifo_store[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15447_ (.CLK(clknet_leaf_81_clk_i),
    .D(_00586_),
    .Q(\fifo0.fifo_store[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15448_ (.CLK(clknet_leaf_85_clk_i),
    .D(_00587_),
    .Q(\fifo0.fifo_store[114][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15449_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00588_),
    .Q(\fifo0.fifo_store[114][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15450_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00589_),
    .Q(\fifo0.fifo_store[114][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15451_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00590_),
    .Q(\fifo0.fifo_store[114][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15452_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00591_),
    .Q(\fifo0.fifo_store[114][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15453_ (.CLK(clknet_leaf_92_clk_i),
    .D(_00592_),
    .Q(\fifo0.fifo_store[114][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15454_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00593_),
    .Q(\fifo0.fifo_store[114][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15455_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00594_),
    .Q(\fifo0.fifo_store[114][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15456_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00595_),
    .Q(\fifo0.fifo_store[114][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15457_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00596_),
    .Q(\fifo0.fifo_store[114][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15458_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00597_),
    .Q(\fifo0.fifo_store[114][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15459_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00598_),
    .Q(\fifo0.fifo_store[114][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15460_ (.CLK(clknet_leaf_56_clk_i),
    .D(_00599_),
    .Q(\fifo0.fifo_store[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15461_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00600_),
    .Q(\fifo0.fifo_store[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15462_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00601_),
    .Q(\fifo0.fifo_store[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15463_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00602_),
    .Q(\fifo0.fifo_store[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15464_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00603_),
    .Q(\fifo0.fifo_store[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15465_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00604_),
    .Q(\fifo0.fifo_store[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15466_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00605_),
    .Q(\fifo0.fifo_store[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15467_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00606_),
    .Q(\fifo0.fifo_store[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15468_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00607_),
    .Q(\fifo0.fifo_store[46][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15469_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00608_),
    .Q(\fifo0.fifo_store[46][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15470_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00609_),
    .Q(\fifo0.fifo_store[46][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15471_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00610_),
    .Q(\fifo0.fifo_store[46][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15472_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00611_),
    .Q(\fifo0.fifo_store[46][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15473_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00612_),
    .Q(\fifo0.fifo_store[46][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15474_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00613_),
    .Q(\fifo0.fifo_store[46][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15475_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00614_),
    .Q(\fifo0.fifo_store[46][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15476_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00615_),
    .Q(\fifo0.fifo_store[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15477_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00616_),
    .Q(\fifo0.fifo_store[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15478_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00617_),
    .Q(\fifo0.fifo_store[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15479_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00618_),
    .Q(\fifo0.fifo_store[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15480_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00619_),
    .Q(\fifo0.fifo_store[91][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15481_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00620_),
    .Q(\fifo0.fifo_store[91][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15482_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00621_),
    .Q(\fifo0.fifo_store[91][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15483_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00622_),
    .Q(\fifo0.fifo_store[91][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15484_ (.CLK(clknet_leaf_134_clk_i),
    .D(_00623_),
    .Q(\fifo0.fifo_store[91][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15485_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00624_),
    .Q(\fifo0.fifo_store[91][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15486_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00625_),
    .Q(\fifo0.fifo_store[91][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15487_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00626_),
    .Q(\fifo0.fifo_store[91][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15488_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00627_),
    .Q(\fifo0.fifo_store[91][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15489_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00628_),
    .Q(\fifo0.fifo_store[91][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15490_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00629_),
    .Q(\fifo0.fifo_store[91][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15491_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00630_),
    .Q(\fifo0.fifo_store[91][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15492_ (.CLK(clknet_leaf_75_clk_i),
    .D(_00631_),
    .Q(\fifo0.fifo_store[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15493_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00632_),
    .Q(\fifo0.fifo_store[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15494_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00633_),
    .Q(\fifo0.fifo_store[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15495_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00634_),
    .Q(\fifo0.fifo_store[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15496_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00635_),
    .Q(\fifo0.fifo_store[66][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15497_ (.CLK(clknet_leaf_103_clk_i),
    .D(_00636_),
    .Q(\fifo0.fifo_store[66][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15498_ (.CLK(clknet_leaf_110_clk_i),
    .D(_00637_),
    .Q(\fifo0.fifo_store[66][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15499_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00638_),
    .Q(\fifo0.fifo_store[66][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15500_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00639_),
    .Q(\fifo0.fifo_store[66][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15501_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00640_),
    .Q(\fifo0.fifo_store[66][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15502_ (.CLK(clknet_leaf_159_clk_i),
    .D(_00641_),
    .Q(\fifo0.fifo_store[66][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15503_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00642_),
    .Q(\fifo0.fifo_store[66][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15504_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00643_),
    .Q(\fifo0.fifo_store[66][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15505_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00644_),
    .Q(\fifo0.fifo_store[66][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15506_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00645_),
    .Q(\fifo0.fifo_store[66][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15507_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00646_),
    .Q(\fifo0.fifo_store[66][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15508_ (.CLK(clknet_leaf_61_clk_i),
    .D(_00647_),
    .Q(\fifo0.fifo_store[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15509_ (.CLK(clknet_leaf_62_clk_i),
    .D(_00648_),
    .Q(\fifo0.fifo_store[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15510_ (.CLK(clknet_leaf_115_clk_i),
    .D(_00649_),
    .Q(\fifo0.fifo_store[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15511_ (.CLK(clknet_leaf_48_clk_i),
    .D(_00650_),
    .Q(\fifo0.fifo_store[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15512_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00651_),
    .Q(\fifo0.fifo_store[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15513_ (.CLK(clknet_leaf_119_clk_i),
    .D(_00652_),
    .Q(\fifo0.fifo_store[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15514_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00653_),
    .Q(\fifo0.fifo_store[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15515_ (.CLK(clknet_leaf_132_clk_i),
    .D(_00654_),
    .Q(\fifo0.fifo_store[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15516_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00655_),
    .Q(\fifo0.fifo_store[49][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15517_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00656_),
    .Q(\fifo0.fifo_store[49][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15518_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00657_),
    .Q(\fifo0.fifo_store[49][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15519_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00658_),
    .Q(\fifo0.fifo_store[49][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15520_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00659_),
    .Q(\fifo0.fifo_store[49][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15521_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00660_),
    .Q(\fifo0.fifo_store[49][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15522_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00661_),
    .Q(\fifo0.fifo_store[49][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15523_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00662_),
    .Q(\fifo0.fifo_store[49][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15524_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00663_),
    .Q(\fifo0.fifo_store[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15525_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00664_),
    .Q(\fifo0.fifo_store[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15526_ (.CLK(clknet_leaf_117_clk_i),
    .D(_00665_),
    .Q(\fifo0.fifo_store[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15527_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00666_),
    .Q(\fifo0.fifo_store[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15528_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00667_),
    .Q(\fifo0.fifo_store[110][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15529_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00668_),
    .Q(\fifo0.fifo_store[110][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15530_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00669_),
    .Q(\fifo0.fifo_store[110][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15531_ (.CLK(clknet_leaf_141_clk_i),
    .D(_00670_),
    .Q(\fifo0.fifo_store[110][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15532_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00671_),
    .Q(\fifo0.fifo_store[110][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15533_ (.CLK(clknet_leaf_113_clk_i),
    .D(_00672_),
    .Q(\fifo0.fifo_store[110][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15534_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00673_),
    .Q(\fifo0.fifo_store[110][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15535_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00674_),
    .Q(\fifo0.fifo_store[110][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15536_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00675_),
    .Q(\fifo0.fifo_store[110][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15537_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00676_),
    .Q(\fifo0.fifo_store[110][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15538_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00677_),
    .Q(\fifo0.fifo_store[110][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15539_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00678_),
    .Q(\fifo0.fifo_store[110][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15540_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00679_),
    .Q(\fifo0.fifo_store[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15541_ (.CLK(clknet_leaf_78_clk_i),
    .D(_00680_),
    .Q(\fifo0.fifo_store[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15542_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00681_),
    .Q(\fifo0.fifo_store[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15543_ (.CLK(clknet_leaf_68_clk_i),
    .D(_00682_),
    .Q(\fifo0.fifo_store[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15544_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00683_),
    .Q(\fifo0.fifo_store[104][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15545_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00684_),
    .Q(\fifo0.fifo_store[104][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15546_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00685_),
    .Q(\fifo0.fifo_store[104][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15547_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00686_),
    .Q(\fifo0.fifo_store[104][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15548_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00687_),
    .Q(\fifo0.fifo_store[104][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15549_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00688_),
    .Q(\fifo0.fifo_store[104][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15550_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00689_),
    .Q(\fifo0.fifo_store[104][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15551_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00690_),
    .Q(\fifo0.fifo_store[104][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15552_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00691_),
    .Q(\fifo0.fifo_store[104][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15553_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00692_),
    .Q(\fifo0.fifo_store[104][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15554_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00693_),
    .Q(\fifo0.fifo_store[104][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15555_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00694_),
    .Q(\fifo0.fifo_store[104][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15556_ (.CLK(clknet_leaf_61_clk_i),
    .D(_00695_),
    .Q(\fifo0.fifo_store[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15557_ (.CLK(clknet_leaf_78_clk_i),
    .D(_00696_),
    .Q(\fifo0.fifo_store[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15558_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00697_),
    .Q(\fifo0.fifo_store[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15559_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00698_),
    .Q(\fifo0.fifo_store[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15560_ (.CLK(clknet_leaf_84_clk_i),
    .D(_00699_),
    .Q(\fifo0.fifo_store[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15561_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00700_),
    .Q(\fifo0.fifo_store[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15562_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00701_),
    .Q(\fifo0.fifo_store[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15563_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00702_),
    .Q(\fifo0.fifo_store[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15564_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00703_),
    .Q(\fifo0.fifo_store[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15565_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00704_),
    .Q(\fifo0.fifo_store[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15566_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00705_),
    .Q(\fifo0.fifo_store[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15567_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00706_),
    .Q(\fifo0.fifo_store[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15568_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00707_),
    .Q(\fifo0.fifo_store[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15569_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00708_),
    .Q(\fifo0.fifo_store[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15570_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00709_),
    .Q(\fifo0.fifo_store[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15571_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00710_),
    .Q(\fifo0.fifo_store[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15572_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00711_),
    .Q(\fifo0.fifo_store[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15573_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00712_),
    .Q(\fifo0.fifo_store[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15574_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00713_),
    .Q(\fifo0.fifo_store[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15575_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00714_),
    .Q(\fifo0.fifo_store[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15576_ (.CLK(clknet_leaf_89_clk_i),
    .D(_00715_),
    .Q(\fifo0.fifo_store[103][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15577_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00716_),
    .Q(\fifo0.fifo_store[103][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15578_ (.CLK(clknet_leaf_110_clk_i),
    .D(_00717_),
    .Q(\fifo0.fifo_store[103][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15579_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00718_),
    .Q(\fifo0.fifo_store[103][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15580_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00719_),
    .Q(\fifo0.fifo_store[103][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15581_ (.CLK(clknet_leaf_45_clk_i),
    .D(_00720_),
    .Q(\fifo0.fifo_store[103][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15582_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00721_),
    .Q(\fifo0.fifo_store[103][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15583_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00722_),
    .Q(\fifo0.fifo_store[103][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15584_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00723_),
    .Q(\fifo0.fifo_store[103][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15585_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00724_),
    .Q(\fifo0.fifo_store[103][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15586_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00725_),
    .Q(\fifo0.fifo_store[103][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15587_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00726_),
    .Q(\fifo0.fifo_store[103][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15588_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00727_),
    .Q(\fifo0.fifo_store[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15589_ (.CLK(clknet_leaf_72_clk_i),
    .D(_00728_),
    .Q(\fifo0.fifo_store[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15590_ (.CLK(clknet_leaf_117_clk_i),
    .D(_00729_),
    .Q(\fifo0.fifo_store[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15591_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00730_),
    .Q(\fifo0.fifo_store[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15592_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00731_),
    .Q(\fifo0.fifo_store[108][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15593_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00732_),
    .Q(\fifo0.fifo_store[108][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15594_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00733_),
    .Q(\fifo0.fifo_store[108][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15595_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00734_),
    .Q(\fifo0.fifo_store[108][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15596_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00735_),
    .Q(\fifo0.fifo_store[108][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15597_ (.CLK(clknet_leaf_88_clk_i),
    .D(_00736_),
    .Q(\fifo0.fifo_store[108][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15598_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00737_),
    .Q(\fifo0.fifo_store[108][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15599_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00738_),
    .Q(\fifo0.fifo_store[108][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15600_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00739_),
    .Q(\fifo0.fifo_store[108][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15601_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00740_),
    .Q(\fifo0.fifo_store[108][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15602_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00741_),
    .Q(\fifo0.fifo_store[108][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15603_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00742_),
    .Q(\fifo0.fifo_store[108][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15604_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00743_),
    .Q(\fifo0.fifo_store[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15605_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00744_),
    .Q(\fifo0.fifo_store[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15606_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00745_),
    .Q(\fifo0.fifo_store[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15607_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00746_),
    .Q(\fifo0.fifo_store[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15608_ (.CLK(clknet_leaf_88_clk_i),
    .D(_00747_),
    .Q(\fifo0.fifo_store[102][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15609_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00748_),
    .Q(\fifo0.fifo_store[102][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15610_ (.CLK(clknet_leaf_111_clk_i),
    .D(_00749_),
    .Q(\fifo0.fifo_store[102][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15611_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00750_),
    .Q(\fifo0.fifo_store[102][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15612_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00751_),
    .Q(\fifo0.fifo_store[102][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15613_ (.CLK(clknet_leaf_113_clk_i),
    .D(_00752_),
    .Q(\fifo0.fifo_store[102][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15614_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00753_),
    .Q(\fifo0.fifo_store[102][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15615_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00754_),
    .Q(\fifo0.fifo_store[102][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15616_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00755_),
    .Q(\fifo0.fifo_store[102][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15617_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00756_),
    .Q(\fifo0.fifo_store[102][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15618_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00757_),
    .Q(\fifo0.fifo_store[102][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15619_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00758_),
    .Q(\fifo0.fifo_store[102][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15620_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00759_),
    .Q(\fifo0.fifo_store[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15621_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00760_),
    .Q(\fifo0.fifo_store[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15622_ (.CLK(clknet_leaf_108_clk_i),
    .D(_00761_),
    .Q(\fifo0.fifo_store[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15623_ (.CLK(clknet_leaf_74_clk_i),
    .D(_00762_),
    .Q(\fifo0.fifo_store[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15624_ (.CLK(clknet_leaf_89_clk_i),
    .D(_00763_),
    .Q(\fifo0.fifo_store[101][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15625_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00764_),
    .Q(\fifo0.fifo_store[101][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15626_ (.CLK(clknet_leaf_111_clk_i),
    .D(_00765_),
    .Q(\fifo0.fifo_store[101][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15627_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00766_),
    .Q(\fifo0.fifo_store[101][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15628_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00767_),
    .Q(\fifo0.fifo_store[101][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15629_ (.CLK(clknet_leaf_114_clk_i),
    .D(_00768_),
    .Q(\fifo0.fifo_store[101][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15630_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00769_),
    .Q(\fifo0.fifo_store[101][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15631_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00770_),
    .Q(\fifo0.fifo_store[101][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15632_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00771_),
    .Q(\fifo0.fifo_store[101][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15633_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00772_),
    .Q(\fifo0.fifo_store[101][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15634_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00773_),
    .Q(\fifo0.fifo_store[101][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15635_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00774_),
    .Q(\fifo0.fifo_store[101][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15636_ (.CLK(clknet_leaf_63_clk_i),
    .D(_00775_),
    .Q(\fifo0.fifo_store[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15637_ (.CLK(clknet_leaf_79_clk_i),
    .D(_00776_),
    .Q(\fifo0.fifo_store[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15638_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00777_),
    .Q(\fifo0.fifo_store[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15639_ (.CLK(clknet_leaf_69_clk_i),
    .D(_00778_),
    .Q(\fifo0.fifo_store[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15640_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00779_),
    .Q(\fifo0.fifo_store[107][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15641_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00780_),
    .Q(\fifo0.fifo_store[107][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15642_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00781_),
    .Q(\fifo0.fifo_store[107][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15643_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00782_),
    .Q(\fifo0.fifo_store[107][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15644_ (.CLK(clknet_leaf_118_clk_i),
    .D(_00783_),
    .Q(\fifo0.fifo_store[107][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15645_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00784_),
    .Q(\fifo0.fifo_store[107][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15646_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00785_),
    .Q(\fifo0.fifo_store[107][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15647_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00786_),
    .Q(\fifo0.fifo_store[107][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15648_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00787_),
    .Q(\fifo0.fifo_store[107][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15649_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00788_),
    .Q(\fifo0.fifo_store[107][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15650_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00789_),
    .Q(\fifo0.fifo_store[107][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15651_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00790_),
    .Q(\fifo0.fifo_store[107][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15652_ (.CLK(clknet_leaf_56_clk_i),
    .D(_00791_),
    .Q(\fifo0.fifo_store[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15653_ (.CLK(clknet_leaf_56_clk_i),
    .D(_00792_),
    .Q(\fifo0.fifo_store[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15654_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00793_),
    .Q(\fifo0.fifo_store[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15655_ (.CLK(clknet_leaf_50_clk_i),
    .D(_00794_),
    .Q(\fifo0.fifo_store[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15656_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00795_),
    .Q(\fifo0.fifo_store[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15657_ (.CLK(clknet_leaf_119_clk_i),
    .D(_00796_),
    .Q(\fifo0.fifo_store[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15658_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00797_),
    .Q(\fifo0.fifo_store[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15659_ (.CLK(clknet_leaf_128_clk_i),
    .D(_00798_),
    .Q(\fifo0.fifo_store[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15660_ (.CLK(clknet_leaf_119_clk_i),
    .D(_00799_),
    .Q(\fifo0.fifo_store[45][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15661_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00800_),
    .Q(\fifo0.fifo_store[45][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15662_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00801_),
    .Q(\fifo0.fifo_store[45][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15663_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00802_),
    .Q(\fifo0.fifo_store[45][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15664_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00803_),
    .Q(\fifo0.fifo_store[45][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15665_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00804_),
    .Q(\fifo0.fifo_store[45][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15666_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00805_),
    .Q(\fifo0.fifo_store[45][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15667_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00806_),
    .Q(\fifo0.fifo_store[45][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15668_ (.CLK(clknet_leaf_72_clk_i),
    .D(_00807_),
    .Q(\fifo0.fifo_store[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15669_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00808_),
    .Q(\fifo0.fifo_store[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15670_ (.CLK(clknet_leaf_109_clk_i),
    .D(_00809_),
    .Q(\fifo0.fifo_store[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15671_ (.CLK(clknet_leaf_69_clk_i),
    .D(_00810_),
    .Q(\fifo0.fifo_store[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15672_ (.CLK(clknet_leaf_88_clk_i),
    .D(_00811_),
    .Q(\fifo0.fifo_store[126][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15673_ (.CLK(clknet_leaf_107_clk_i),
    .D(_00812_),
    .Q(\fifo0.fifo_store[126][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15674_ (.CLK(clknet_leaf_111_clk_i),
    .D(_00813_),
    .Q(\fifo0.fifo_store[126][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15675_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00814_),
    .Q(\fifo0.fifo_store[126][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15676_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00815_),
    .Q(\fifo0.fifo_store[126][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15677_ (.CLK(clknet_leaf_88_clk_i),
    .D(_00816_),
    .Q(\fifo0.fifo_store[126][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15678_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00817_),
    .Q(\fifo0.fifo_store[126][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15679_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00818_),
    .Q(\fifo0.fifo_store[126][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15680_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00819_),
    .Q(\fifo0.fifo_store[126][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15681_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00820_),
    .Q(\fifo0.fifo_store[126][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15682_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00821_),
    .Q(\fifo0.fifo_store[126][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15683_ (.CLK(clknet_leaf_157_clk_i),
    .D(_00822_),
    .Q(\fifo0.fifo_store[126][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15684_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00823_),
    .Q(\fifo0.fifo_store[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15685_ (.CLK(clknet_leaf_71_clk_i),
    .D(_00824_),
    .Q(\fifo0.fifo_store[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15686_ (.CLK(clknet_leaf_109_clk_i),
    .D(_00825_),
    .Q(\fifo0.fifo_store[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15687_ (.CLK(clknet_leaf_68_clk_i),
    .D(_00826_),
    .Q(\fifo0.fifo_store[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15688_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00827_),
    .Q(\fifo0.fifo_store[125][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15689_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00828_),
    .Q(\fifo0.fifo_store[125][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15690_ (.CLK(clknet_leaf_112_clk_i),
    .D(_00829_),
    .Q(\fifo0.fifo_store[125][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15691_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00830_),
    .Q(\fifo0.fifo_store[125][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15692_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00831_),
    .Q(\fifo0.fifo_store[125][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15693_ (.CLK(clknet_leaf_89_clk_i),
    .D(_00832_),
    .Q(\fifo0.fifo_store[125][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15694_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00833_),
    .Q(\fifo0.fifo_store[125][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15695_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00834_),
    .Q(\fifo0.fifo_store[125][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15696_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00835_),
    .Q(\fifo0.fifo_store[125][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15697_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00836_),
    .Q(\fifo0.fifo_store[125][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15698_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00837_),
    .Q(\fifo0.fifo_store[125][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15699_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00838_),
    .Q(\fifo0.fifo_store[125][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15700_ (.CLK(clknet_leaf_75_clk_i),
    .D(_00839_),
    .Q(\fifo0.fifo_store[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15701_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00840_),
    .Q(\fifo0.fifo_store[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15702_ (.CLK(clknet_leaf_106_clk_i),
    .D(_00841_),
    .Q(\fifo0.fifo_store[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15703_ (.CLK(clknet_leaf_77_clk_i),
    .D(_00842_),
    .Q(\fifo0.fifo_store[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15704_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00843_),
    .Q(\fifo0.fifo_store[65][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15705_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00844_),
    .Q(\fifo0.fifo_store[65][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15706_ (.CLK(clknet_leaf_110_clk_i),
    .D(_00845_),
    .Q(\fifo0.fifo_store[65][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15707_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00846_),
    .Q(\fifo0.fifo_store[65][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15708_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00847_),
    .Q(\fifo0.fifo_store[65][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15709_ (.CLK(clknet_leaf_90_clk_i),
    .D(_00848_),
    .Q(\fifo0.fifo_store[65][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15710_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00849_),
    .Q(\fifo0.fifo_store[65][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15711_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00850_),
    .Q(\fifo0.fifo_store[65][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15712_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00851_),
    .Q(\fifo0.fifo_store[65][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15713_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00852_),
    .Q(\fifo0.fifo_store[65][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15714_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00853_),
    .Q(\fifo0.fifo_store[65][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15715_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00854_),
    .Q(\fifo0.fifo_store[65][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15716_ (.CLK(clknet_leaf_75_clk_i),
    .D(_00855_),
    .Q(\fifo0.fifo_store[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15717_ (.CLK(clknet_leaf_76_clk_i),
    .D(_00856_),
    .Q(\fifo0.fifo_store[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15718_ (.CLK(clknet_leaf_103_clk_i),
    .D(_00857_),
    .Q(\fifo0.fifo_store[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15719_ (.CLK(clknet_leaf_77_clk_i),
    .D(_00858_),
    .Q(\fifo0.fifo_store[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15720_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00859_),
    .Q(\fifo0.fifo_store[64][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15721_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00860_),
    .Q(\fifo0.fifo_store[64][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15722_ (.CLK(clknet_leaf_105_clk_i),
    .D(_00861_),
    .Q(\fifo0.fifo_store[64][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15723_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00862_),
    .Q(\fifo0.fifo_store[64][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15724_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00863_),
    .Q(\fifo0.fifo_store[64][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15725_ (.CLK(clknet_leaf_89_clk_i),
    .D(_00864_),
    .Q(\fifo0.fifo_store[64][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15726_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00865_),
    .Q(\fifo0.fifo_store[64][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15727_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00866_),
    .Q(\fifo0.fifo_store[64][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15728_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00867_),
    .Q(\fifo0.fifo_store[64][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15729_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00868_),
    .Q(\fifo0.fifo_store[64][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15730_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00869_),
    .Q(\fifo0.fifo_store[64][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15731_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00870_),
    .Q(\fifo0.fifo_store[64][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15732_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00871_),
    .Q(\fifo0.fifo_store[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15733_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00872_),
    .Q(\fifo0.fifo_store[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15734_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00873_),
    .Q(\fifo0.fifo_store[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15735_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00874_),
    .Q(\fifo0.fifo_store[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15736_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00875_),
    .Q(\fifo0.fifo_store[90][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15737_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00876_),
    .Q(\fifo0.fifo_store[90][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15738_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00877_),
    .Q(\fifo0.fifo_store[90][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15739_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00878_),
    .Q(\fifo0.fifo_store[90][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15740_ (.CLK(clknet_leaf_134_clk_i),
    .D(_00879_),
    .Q(\fifo0.fifo_store[90][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15741_ (.CLK(clknet_leaf_45_clk_i),
    .D(_00880_),
    .Q(\fifo0.fifo_store[90][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15742_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00881_),
    .Q(\fifo0.fifo_store[90][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15743_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00882_),
    .Q(\fifo0.fifo_store[90][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15744_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00883_),
    .Q(\fifo0.fifo_store[90][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15745_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00884_),
    .Q(\fifo0.fifo_store[90][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15746_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00885_),
    .Q(\fifo0.fifo_store[90][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15747_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00886_),
    .Q(\fifo0.fifo_store[90][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15748_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00887_),
    .Q(\fifo0.fifo_store[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15749_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00888_),
    .Q(\fifo0.fifo_store[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15750_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00889_),
    .Q(\fifo0.fifo_store[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15751_ (.CLK(clknet_leaf_66_clk_i),
    .D(_00890_),
    .Q(\fifo0.fifo_store[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15752_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00891_),
    .Q(\fifo0.fifo_store[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15753_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00892_),
    .Q(\fifo0.fifo_store[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15754_ (.CLK(clknet_leaf_102_clk_i),
    .D(_00893_),
    .Q(\fifo0.fifo_store[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15755_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00894_),
    .Q(\fifo0.fifo_store[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15756_ (.CLK(clknet_leaf_126_clk_i),
    .D(_00895_),
    .Q(\fifo0.fifo_store[63][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15757_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00896_),
    .Q(\fifo0.fifo_store[63][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15758_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00897_),
    .Q(\fifo0.fifo_store[63][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15759_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00898_),
    .Q(\fifo0.fifo_store[63][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15760_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00899_),
    .Q(\fifo0.fifo_store[63][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15761_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00900_),
    .Q(\fifo0.fifo_store[63][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15762_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00901_),
    .Q(\fifo0.fifo_store[63][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15763_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00902_),
    .Q(\fifo0.fifo_store[63][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15764_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00903_),
    .Q(\fifo0.fifo_store[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15765_ (.CLK(clknet_leaf_55_clk_i),
    .D(_00904_),
    .Q(\fifo0.fifo_store[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15766_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00905_),
    .Q(\fifo0.fifo_store[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15767_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00906_),
    .Q(\fifo0.fifo_store[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15768_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00907_),
    .Q(\fifo0.fifo_store[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15769_ (.CLK(clknet_leaf_101_clk_i),
    .D(_00908_),
    .Q(\fifo0.fifo_store[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15770_ (.CLK(clknet_leaf_103_clk_i),
    .D(_00909_),
    .Q(\fifo0.fifo_store[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15771_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00910_),
    .Q(\fifo0.fifo_store[62][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15772_ (.CLK(clknet_leaf_119_clk_i),
    .D(_00911_),
    .Q(\fifo0.fifo_store[62][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15773_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00912_),
    .Q(\fifo0.fifo_store[62][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15774_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00913_),
    .Q(\fifo0.fifo_store[62][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15775_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00914_),
    .Q(\fifo0.fifo_store[62][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15776_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00915_),
    .Q(\fifo0.fifo_store[62][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15777_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00916_),
    .Q(\fifo0.fifo_store[62][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15778_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00917_),
    .Q(\fifo0.fifo_store[62][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15779_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00918_),
    .Q(\fifo0.fifo_store[62][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15780_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00919_),
    .Q(\fifo0.fifo_store[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15781_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00920_),
    .Q(\fifo0.fifo_store[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15782_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00921_),
    .Q(\fifo0.fifo_store[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15783_ (.CLK(clknet_leaf_87_clk_i),
    .D(_00922_),
    .Q(\fifo0.fifo_store[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15784_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00923_),
    .Q(\fifo0.fifo_store[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15785_ (.CLK(clknet_leaf_146_clk_i),
    .D(_00924_),
    .Q(\fifo0.fifo_store[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15786_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00925_),
    .Q(\fifo0.fifo_store[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15787_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00926_),
    .Q(\fifo0.fifo_store[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15788_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00927_),
    .Q(\fifo0.fifo_store[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15789_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00928_),
    .Q(\fifo0.fifo_store[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15790_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00929_),
    .Q(\fifo0.fifo_store[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15791_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00930_),
    .Q(\fifo0.fifo_store[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15792_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00931_),
    .Q(\fifo0.fifo_store[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15793_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00932_),
    .Q(\fifo0.fifo_store[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15794_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00933_),
    .Q(\fifo0.fifo_store[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15795_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00934_),
    .Q(\fifo0.fifo_store[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15796_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00935_),
    .Q(\fifo0.fifo_store[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15797_ (.CLK(clknet_leaf_49_clk_i),
    .D(_00936_),
    .Q(\fifo0.fifo_store[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15798_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00937_),
    .Q(\fifo0.fifo_store[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15799_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00938_),
    .Q(\fifo0.fifo_store[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15800_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00939_),
    .Q(\fifo0.fifo_store[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15801_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00940_),
    .Q(\fifo0.fifo_store[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15802_ (.CLK(clknet_leaf_102_clk_i),
    .D(_00941_),
    .Q(\fifo0.fifo_store[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15803_ (.CLK(clknet_leaf_149_clk_i),
    .D(_00942_),
    .Q(\fifo0.fifo_store[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15804_ (.CLK(clknet_leaf_122_clk_i),
    .D(_00943_),
    .Q(\fifo0.fifo_store[61][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15805_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00944_),
    .Q(\fifo0.fifo_store[61][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15806_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00945_),
    .Q(\fifo0.fifo_store[61][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15807_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00946_),
    .Q(\fifo0.fifo_store[61][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15808_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00947_),
    .Q(\fifo0.fifo_store[61][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15809_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00948_),
    .Q(\fifo0.fifo_store[61][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15810_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00949_),
    .Q(\fifo0.fifo_store[61][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15811_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00950_),
    .Q(\fifo0.fifo_store[61][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15812_ (.CLK(clknet_leaf_65_clk_i),
    .D(_00951_),
    .Q(\fifo0.fifo_store[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15813_ (.CLK(clknet_leaf_49_clk_i),
    .D(_00952_),
    .Q(\fifo0.fifo_store[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15814_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00953_),
    .Q(\fifo0.fifo_store[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15815_ (.CLK(clknet_leaf_46_clk_i),
    .D(_00954_),
    .Q(\fifo0.fifo_store[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15816_ (.CLK(clknet_leaf_94_clk_i),
    .D(_00955_),
    .Q(\fifo0.fifo_store[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15817_ (.CLK(clknet_leaf_148_clk_i),
    .D(_00956_),
    .Q(\fifo0.fifo_store[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15818_ (.CLK(clknet_leaf_102_clk_i),
    .D(_00957_),
    .Q(\fifo0.fifo_store[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15819_ (.CLK(clknet_leaf_149_clk_i),
    .D(_00958_),
    .Q(\fifo0.fifo_store[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15820_ (.CLK(clknet_leaf_119_clk_i),
    .D(_00959_),
    .Q(\fifo0.fifo_store[60][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15821_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00960_),
    .Q(\fifo0.fifo_store[60][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15822_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00961_),
    .Q(\fifo0.fifo_store[60][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15823_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00962_),
    .Q(\fifo0.fifo_store[60][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15824_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00963_),
    .Q(\fifo0.fifo_store[60][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15825_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00964_),
    .Q(\fifo0.fifo_store[60][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15826_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00965_),
    .Q(\fifo0.fifo_store[60][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15827_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00966_),
    .Q(\fifo0.fifo_store[60][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15828_ (.CLK(clknet_leaf_64_clk_i),
    .D(_00967_),
    .Q(\fifo0.fifo_store[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15829_ (.CLK(clknet_leaf_80_clk_i),
    .D(_00968_),
    .Q(\fifo0.fifo_store[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15830_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00969_),
    .Q(\fifo0.fifo_store[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15831_ (.CLK(clknet_leaf_86_clk_i),
    .D(_00970_),
    .Q(\fifo0.fifo_store[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15832_ (.CLK(clknet_leaf_93_clk_i),
    .D(_00971_),
    .Q(\fifo0.fifo_store[88][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15833_ (.CLK(clknet_leaf_147_clk_i),
    .D(_00972_),
    .Q(\fifo0.fifo_store[88][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15834_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00973_),
    .Q(\fifo0.fifo_store[88][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15835_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00974_),
    .Q(\fifo0.fifo_store[88][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15836_ (.CLK(clknet_leaf_133_clk_i),
    .D(_00975_),
    .Q(\fifo0.fifo_store[88][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15837_ (.CLK(clknet_leaf_43_clk_i),
    .D(_00976_),
    .Q(\fifo0.fifo_store[88][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15838_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00977_),
    .Q(\fifo0.fifo_store[88][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15839_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00978_),
    .Q(\fifo0.fifo_store[88][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15840_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00979_),
    .Q(\fifo0.fifo_store[88][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15841_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00980_),
    .Q(\fifo0.fifo_store[88][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15842_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00981_),
    .Q(\fifo0.fifo_store[88][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15843_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00982_),
    .Q(\fifo0.fifo_store[88][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15844_ (.CLK(clknet_leaf_53_clk_i),
    .D(_00983_),
    .Q(\fifo0.fifo_store[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15845_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00984_),
    .Q(\fifo0.fifo_store[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15846_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00985_),
    .Q(\fifo0.fifo_store[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15847_ (.CLK(clknet_leaf_52_clk_i),
    .D(_00986_),
    .Q(\fifo0.fifo_store[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15848_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00987_),
    .Q(\fifo0.fifo_store[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15849_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00988_),
    .Q(\fifo0.fifo_store[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15850_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00989_),
    .Q(\fifo0.fifo_store[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15851_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00990_),
    .Q(\fifo0.fifo_store[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15852_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00991_),
    .Q(\fifo0.fifo_store[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15853_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00992_),
    .Q(\fifo0.fifo_store[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15854_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00993_),
    .Q(\fifo0.fifo_store[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15855_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00994_),
    .Q(\fifo0.fifo_store[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15856_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00995_),
    .Q(\fifo0.fifo_store[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15857_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00996_),
    .Q(\fifo0.fifo_store[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15858_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00997_),
    .Q(\fifo0.fifo_store[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15859_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00998_),
    .Q(\fifo0.fifo_store[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15860_ (.CLK(clknet_leaf_53_clk_i),
    .D(_00999_),
    .Q(\fifo0.fifo_store[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15861_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01000_),
    .Q(\fifo0.fifo_store[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15862_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01001_),
    .Q(\fifo0.fifo_store[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15863_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01002_),
    .Q(\fifo0.fifo_store[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15864_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01003_),
    .Q(\fifo0.fifo_store[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15865_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01004_),
    .Q(\fifo0.fifo_store[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15866_ (.CLK(clknet_leaf_33_clk_i),
    .D(_01005_),
    .Q(\fifo0.fifo_store[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15867_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01006_),
    .Q(\fifo0.fifo_store[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15868_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01007_),
    .Q(\fifo0.fifo_store[58][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15869_ (.CLK(clknet_leaf_39_clk_i),
    .D(_01008_),
    .Q(\fifo0.fifo_store[58][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15870_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01009_),
    .Q(\fifo0.fifo_store[58][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15871_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01010_),
    .Q(\fifo0.fifo_store[58][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15872_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01011_),
    .Q(\fifo0.fifo_store[58][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15873_ (.CLK(clknet_leaf_235_clk_i),
    .D(_01012_),
    .Q(\fifo0.fifo_store[58][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15874_ (.CLK(clknet_leaf_235_clk_i),
    .D(_01013_),
    .Q(\fifo0.fifo_store[58][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15875_ (.CLK(clknet_leaf_219_clk_i),
    .D(_01014_),
    .Q(\fifo0.fifo_store[58][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15876_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01015_),
    .Q(\fifo0.fifo_store[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15877_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01016_),
    .Q(\fifo0.fifo_store[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15878_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01017_),
    .Q(\fifo0.fifo_store[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15879_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01018_),
    .Q(\fifo0.fifo_store[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15880_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01019_),
    .Q(\fifo0.fifo_store[87][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15881_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01020_),
    .Q(\fifo0.fifo_store[87][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15882_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01021_),
    .Q(\fifo0.fifo_store[87][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15883_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01022_),
    .Q(\fifo0.fifo_store[87][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15884_ (.CLK(clknet_leaf_212_clk_i),
    .D(_01023_),
    .Q(\fifo0.fifo_store[87][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15885_ (.CLK(clknet_leaf_42_clk_i),
    .D(_01024_),
    .Q(\fifo0.fifo_store[87][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15886_ (.CLK(clknet_leaf_209_clk_i),
    .D(_01025_),
    .Q(\fifo0.fifo_store[87][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15887_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01026_),
    .Q(\fifo0.fifo_store[87][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15888_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01027_),
    .Q(\fifo0.fifo_store[87][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15889_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01028_),
    .Q(\fifo0.fifo_store[87][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15890_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01029_),
    .Q(\fifo0.fifo_store[87][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15891_ (.CLK(clknet_leaf_211_clk_i),
    .D(_01030_),
    .Q(\fifo0.fifo_store[87][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15892_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01031_),
    .Q(\fifo0.fifo_store[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15893_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01032_),
    .Q(\fifo0.fifo_store[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15894_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01033_),
    .Q(\fifo0.fifo_store[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15895_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01034_),
    .Q(\fifo0.fifo_store[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15896_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01035_),
    .Q(\fifo0.fifo_store[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15897_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01036_),
    .Q(\fifo0.fifo_store[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15898_ (.CLK(clknet_leaf_33_clk_i),
    .D(_01037_),
    .Q(\fifo0.fifo_store[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15899_ (.CLK(clknet_leaf_132_clk_i),
    .D(_01038_),
    .Q(\fifo0.fifo_store[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15900_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01039_),
    .Q(\fifo0.fifo_store[57][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15901_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01040_),
    .Q(\fifo0.fifo_store[57][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15902_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01041_),
    .Q(\fifo0.fifo_store[57][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15903_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01042_),
    .Q(\fifo0.fifo_store[57][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15904_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01043_),
    .Q(\fifo0.fifo_store[57][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15905_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01044_),
    .Q(\fifo0.fifo_store[57][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15906_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01045_),
    .Q(\fifo0.fifo_store[57][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15907_ (.CLK(clknet_leaf_221_clk_i),
    .D(_01046_),
    .Q(\fifo0.fifo_store[57][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15908_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01047_),
    .Q(\fifo0.fifo_store[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15909_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01048_),
    .Q(\fifo0.fifo_store[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15910_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01049_),
    .Q(\fifo0.fifo_store[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15911_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01050_),
    .Q(\fifo0.fifo_store[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15912_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01051_),
    .Q(\fifo0.fifo_store[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15913_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01052_),
    .Q(\fifo0.fifo_store[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15914_ (.CLK(clknet_leaf_33_clk_i),
    .D(_01053_),
    .Q(\fifo0.fifo_store[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15915_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01054_),
    .Q(\fifo0.fifo_store[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15916_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01055_),
    .Q(\fifo0.fifo_store[56][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15917_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01056_),
    .Q(\fifo0.fifo_store[56][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15918_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01057_),
    .Q(\fifo0.fifo_store[56][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15919_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01058_),
    .Q(\fifo0.fifo_store[56][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15920_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01059_),
    .Q(\fifo0.fifo_store[56][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15921_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01060_),
    .Q(\fifo0.fifo_store[56][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15922_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01061_),
    .Q(\fifo0.fifo_store[56][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15923_ (.CLK(clknet_leaf_221_clk_i),
    .D(_01062_),
    .Q(\fifo0.fifo_store[56][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15924_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01063_),
    .Q(\fifo0.fifo_store[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15925_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01064_),
    .Q(\fifo0.fifo_store[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15926_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01065_),
    .Q(\fifo0.fifo_store[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15927_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01066_),
    .Q(\fifo0.fifo_store[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15928_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01067_),
    .Q(\fifo0.fifo_store[86][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15929_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01068_),
    .Q(\fifo0.fifo_store[86][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15930_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01069_),
    .Q(\fifo0.fifo_store[86][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15931_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01070_),
    .Q(\fifo0.fifo_store[86][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15932_ (.CLK(clknet_leaf_212_clk_i),
    .D(_01071_),
    .Q(\fifo0.fifo_store[86][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15933_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01072_),
    .Q(\fifo0.fifo_store[86][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15934_ (.CLK(clknet_leaf_209_clk_i),
    .D(_01073_),
    .Q(\fifo0.fifo_store[86][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15935_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01074_),
    .Q(\fifo0.fifo_store[86][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15936_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01075_),
    .Q(\fifo0.fifo_store[86][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15937_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01076_),
    .Q(\fifo0.fifo_store[86][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15938_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01077_),
    .Q(\fifo0.fifo_store[86][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15939_ (.CLK(clknet_leaf_211_clk_i),
    .D(_01078_),
    .Q(\fifo0.fifo_store[86][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15940_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01079_),
    .Q(\fifo0.fifo_store[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15941_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01080_),
    .Q(\fifo0.fifo_store[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15942_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01081_),
    .Q(\fifo0.fifo_store[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15943_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01082_),
    .Q(\fifo0.fifo_store[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15944_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01083_),
    .Q(\fifo0.fifo_store[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15945_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01084_),
    .Q(\fifo0.fifo_store[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15946_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01085_),
    .Q(\fifo0.fifo_store[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15947_ (.CLK(clknet_leaf_151_clk_i),
    .D(_01086_),
    .Q(\fifo0.fifo_store[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15948_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01087_),
    .Q(\fifo0.fifo_store[55][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15949_ (.CLK(clknet_leaf_37_clk_i),
    .D(_01088_),
    .Q(\fifo0.fifo_store[55][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15950_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01089_),
    .Q(\fifo0.fifo_store[55][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15951_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01090_),
    .Q(\fifo0.fifo_store[55][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15952_ (.CLK(clknet_leaf_234_clk_i),
    .D(_01091_),
    .Q(\fifo0.fifo_store[55][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15953_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01092_),
    .Q(\fifo0.fifo_store[55][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15954_ (.CLK(clknet_leaf_234_clk_i),
    .D(_01093_),
    .Q(\fifo0.fifo_store[55][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15955_ (.CLK(clknet_leaf_221_clk_i),
    .D(_01094_),
    .Q(\fifo0.fifo_store[55][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15956_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01095_),
    .Q(\fifo0.fifo_store[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15957_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01096_),
    .Q(\fifo0.fifo_store[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15958_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01097_),
    .Q(\fifo0.fifo_store[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15959_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01098_),
    .Q(\fifo0.fifo_store[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15960_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01099_),
    .Q(\fifo0.fifo_store[85][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15961_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01100_),
    .Q(\fifo0.fifo_store[85][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15962_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01101_),
    .Q(\fifo0.fifo_store[85][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15963_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01102_),
    .Q(\fifo0.fifo_store[85][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15964_ (.CLK(clknet_leaf_213_clk_i),
    .D(_01103_),
    .Q(\fifo0.fifo_store[85][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15965_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01104_),
    .Q(\fifo0.fifo_store[85][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15966_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01105_),
    .Q(\fifo0.fifo_store[85][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15967_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01106_),
    .Q(\fifo0.fifo_store[85][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15968_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01107_),
    .Q(\fifo0.fifo_store[85][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15969_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01108_),
    .Q(\fifo0.fifo_store[85][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15970_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01109_),
    .Q(\fifo0.fifo_store[85][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15971_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01110_),
    .Q(\fifo0.fifo_store[85][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15972_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01111_),
    .Q(\fifo0.fifo_store[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15973_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01112_),
    .Q(\fifo0.fifo_store[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15974_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01113_),
    .Q(\fifo0.fifo_store[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15975_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01114_),
    .Q(\fifo0.fifo_store[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15976_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01115_),
    .Q(\fifo0.fifo_store[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15977_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01116_),
    .Q(\fifo0.fifo_store[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15978_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01117_),
    .Q(\fifo0.fifo_store[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15979_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01118_),
    .Q(\fifo0.fifo_store[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15980_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01119_),
    .Q(\fifo0.fifo_store[54][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15981_ (.CLK(clknet_leaf_37_clk_i),
    .D(_01120_),
    .Q(\fifo0.fifo_store[54][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15982_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01121_),
    .Q(\fifo0.fifo_store[54][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15983_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01122_),
    .Q(\fifo0.fifo_store[54][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15984_ (.CLK(clknet_leaf_235_clk_i),
    .D(_01123_),
    .Q(\fifo0.fifo_store[54][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15985_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01124_),
    .Q(\fifo0.fifo_store[54][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15986_ (.CLK(clknet_leaf_235_clk_i),
    .D(_01125_),
    .Q(\fifo0.fifo_store[54][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15987_ (.CLK(clknet_leaf_211_clk_i),
    .D(_01126_),
    .Q(\fifo0.fifo_store[54][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15988_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01127_),
    .Q(\fifo0.fifo_store[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15989_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01128_),
    .Q(\fifo0.fifo_store[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15990_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01129_),
    .Q(\fifo0.fifo_store[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15991_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01130_),
    .Q(\fifo0.fifo_store[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15992_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01131_),
    .Q(\fifo0.fifo_store[84][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15993_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01132_),
    .Q(\fifo0.fifo_store[84][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15994_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01133_),
    .Q(\fifo0.fifo_store[84][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15995_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01134_),
    .Q(\fifo0.fifo_store[84][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15996_ (.CLK(clknet_leaf_213_clk_i),
    .D(_01135_),
    .Q(\fifo0.fifo_store[84][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15997_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01136_),
    .Q(\fifo0.fifo_store[84][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15998_ (.CLK(clknet_leaf_209_clk_i),
    .D(_01137_),
    .Q(\fifo0.fifo_store[84][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15999_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01138_),
    .Q(\fifo0.fifo_store[84][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16000_ (.CLK(clknet_leaf_189_clk_i),
    .D(_01139_),
    .Q(\fifo0.fifo_store[84][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16001_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01140_),
    .Q(\fifo0.fifo_store[84][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16002_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01141_),
    .Q(\fifo0.fifo_store[84][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16003_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01142_),
    .Q(\fifo0.fifo_store[84][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16004_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01143_),
    .Q(\fifo0.fifo_store[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16005_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01144_),
    .Q(\fifo0.fifo_store[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16006_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01145_),
    .Q(\fifo0.fifo_store[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16007_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01146_),
    .Q(\fifo0.fifo_store[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16008_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01147_),
    .Q(\fifo0.fifo_store[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16009_ (.CLK(clknet_leaf_207_clk_i),
    .D(_01148_),
    .Q(\fifo0.fifo_store[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16010_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01149_),
    .Q(\fifo0.fifo_store[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16011_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01150_),
    .Q(\fifo0.fifo_store[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16012_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01151_),
    .Q(\fifo0.fifo_store[53][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16013_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01152_),
    .Q(\fifo0.fifo_store[53][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16014_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01153_),
    .Q(\fifo0.fifo_store[53][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16015_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01154_),
    .Q(\fifo0.fifo_store[53][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16016_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01155_),
    .Q(\fifo0.fifo_store[53][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16017_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01156_),
    .Q(\fifo0.fifo_store[53][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16018_ (.CLK(clknet_leaf_232_clk_i),
    .D(_01157_),
    .Q(\fifo0.fifo_store[53][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16019_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01158_),
    .Q(\fifo0.fifo_store[53][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16020_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01159_),
    .Q(\fifo0.fifo_store[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16021_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01160_),
    .Q(\fifo0.fifo_store[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16022_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01161_),
    .Q(\fifo0.fifo_store[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16023_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01162_),
    .Q(\fifo0.fifo_store[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16024_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01163_),
    .Q(\fifo0.fifo_store[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16025_ (.CLK(clknet_leaf_207_clk_i),
    .D(_01164_),
    .Q(\fifo0.fifo_store[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16026_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01165_),
    .Q(\fifo0.fifo_store[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16027_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01166_),
    .Q(\fifo0.fifo_store[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16028_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01167_),
    .Q(\fifo0.fifo_store[52][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16029_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01168_),
    .Q(\fifo0.fifo_store[52][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16030_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01169_),
    .Q(\fifo0.fifo_store[52][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16031_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01170_),
    .Q(\fifo0.fifo_store[52][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16032_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01171_),
    .Q(\fifo0.fifo_store[52][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16033_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01172_),
    .Q(\fifo0.fifo_store[52][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16034_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01173_),
    .Q(\fifo0.fifo_store[52][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16035_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01174_),
    .Q(\fifo0.fifo_store[52][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16036_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01175_),
    .Q(\fifo0.fifo_store[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16037_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01176_),
    .Q(\fifo0.fifo_store[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16038_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01177_),
    .Q(\fifo0.fifo_store[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16039_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01178_),
    .Q(\fifo0.fifo_store[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16040_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01179_),
    .Q(\fifo0.fifo_store[83][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16041_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01180_),
    .Q(\fifo0.fifo_store[83][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16042_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01181_),
    .Q(\fifo0.fifo_store[83][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16043_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01182_),
    .Q(\fifo0.fifo_store[83][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16044_ (.CLK(clknet_leaf_214_clk_i),
    .D(_01183_),
    .Q(\fifo0.fifo_store[83][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16045_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01184_),
    .Q(\fifo0.fifo_store[83][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16046_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01185_),
    .Q(\fifo0.fifo_store[83][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16047_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01186_),
    .Q(\fifo0.fifo_store[83][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16048_ (.CLK(clknet_leaf_238_clk_i),
    .D(_01187_),
    .Q(\fifo0.fifo_store[83][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16049_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01188_),
    .Q(\fifo0.fifo_store[83][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16050_ (.CLK(clknet_leaf_238_clk_i),
    .D(_01189_),
    .Q(\fifo0.fifo_store[83][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16051_ (.CLK(clknet_leaf_211_clk_i),
    .D(_01190_),
    .Q(\fifo0.fifo_store[83][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16052_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01191_),
    .Q(\fifo0.fifo_store[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16053_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01192_),
    .Q(\fifo0.fifo_store[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16054_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01193_),
    .Q(\fifo0.fifo_store[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16055_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01194_),
    .Q(\fifo0.fifo_store[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16056_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01195_),
    .Q(\fifo0.fifo_store[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16057_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01196_),
    .Q(\fifo0.fifo_store[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16058_ (.CLK(clknet_leaf_35_clk_i),
    .D(_01197_),
    .Q(\fifo0.fifo_store[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16059_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01198_),
    .Q(\fifo0.fifo_store[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16060_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01199_),
    .Q(\fifo0.fifo_store[51][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16061_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01200_),
    .Q(\fifo0.fifo_store[51][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16062_ (.CLK(clknet_leaf_222_clk_i),
    .D(_01201_),
    .Q(\fifo0.fifo_store[51][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16063_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01202_),
    .Q(\fifo0.fifo_store[51][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16064_ (.CLK(clknet_leaf_231_clk_i),
    .D(_01203_),
    .Q(\fifo0.fifo_store[51][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16065_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01204_),
    .Q(\fifo0.fifo_store[51][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16066_ (.CLK(clknet_leaf_234_clk_i),
    .D(_01205_),
    .Q(\fifo0.fifo_store[51][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16067_ (.CLK(clknet_leaf_221_clk_i),
    .D(_01206_),
    .Q(\fifo0.fifo_store[51][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16068_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01207_),
    .Q(\fifo0.fifo_store[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16069_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01208_),
    .Q(\fifo0.fifo_store[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16070_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01209_),
    .Q(\fifo0.fifo_store[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16071_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01210_),
    .Q(\fifo0.fifo_store[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16072_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01211_),
    .Q(\fifo0.fifo_store[106][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16073_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01212_),
    .Q(\fifo0.fifo_store[106][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16074_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01213_),
    .Q(\fifo0.fifo_store[106][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16075_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01214_),
    .Q(\fifo0.fifo_store[106][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16076_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01215_),
    .Q(\fifo0.fifo_store[106][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16077_ (.CLK(clknet_leaf_44_clk_i),
    .D(_01216_),
    .Q(\fifo0.fifo_store[106][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16078_ (.CLK(clknet_leaf_197_clk_i),
    .D(_01217_),
    .Q(\fifo0.fifo_store[106][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16079_ (.CLK(clknet_leaf_180_clk_i),
    .D(_01218_),
    .Q(\fifo0.fifo_store[106][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16080_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01219_),
    .Q(\fifo0.fifo_store[106][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16081_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01220_),
    .Q(\fifo0.fifo_store[106][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16082_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01221_),
    .Q(\fifo0.fifo_store[106][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16083_ (.CLK(clknet_leaf_134_clk_i),
    .D(_01222_),
    .Q(\fifo0.fifo_store[106][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16084_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01223_),
    .Q(\fifo0.fifo_store[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16085_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01224_),
    .Q(\fifo0.fifo_store[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16086_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01225_),
    .Q(\fifo0.fifo_store[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16087_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01226_),
    .Q(\fifo0.fifo_store[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16088_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01227_),
    .Q(\fifo0.fifo_store[82][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16089_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01228_),
    .Q(\fifo0.fifo_store[82][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16090_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01229_),
    .Q(\fifo0.fifo_store[82][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16091_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01230_),
    .Q(\fifo0.fifo_store[82][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16092_ (.CLK(clknet_leaf_214_clk_i),
    .D(_01231_),
    .Q(\fifo0.fifo_store[82][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16093_ (.CLK(clknet_leaf_42_clk_i),
    .D(_01232_),
    .Q(\fifo0.fifo_store[82][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16094_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01233_),
    .Q(\fifo0.fifo_store[82][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16095_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01234_),
    .Q(\fifo0.fifo_store[82][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16096_ (.CLK(clknet_leaf_239_clk_i),
    .D(_01235_),
    .Q(\fifo0.fifo_store[82][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16097_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01236_),
    .Q(\fifo0.fifo_store[82][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16098_ (.CLK(clknet_leaf_238_clk_i),
    .D(_01237_),
    .Q(\fifo0.fifo_store[82][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16099_ (.CLK(clknet_leaf_214_clk_i),
    .D(_01238_),
    .Q(\fifo0.fifo_store[82][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16100_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01239_),
    .Q(\fifo0.fifo_store[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16101_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01240_),
    .Q(\fifo0.fifo_store[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16102_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01241_),
    .Q(\fifo0.fifo_store[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16103_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01242_),
    .Q(\fifo0.fifo_store[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16104_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01243_),
    .Q(\fifo0.fifo_store[81][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16105_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01244_),
    .Q(\fifo0.fifo_store[81][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16106_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01245_),
    .Q(\fifo0.fifo_store[81][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16107_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01246_),
    .Q(\fifo0.fifo_store[81][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16108_ (.CLK(clknet_leaf_213_clk_i),
    .D(_01247_),
    .Q(\fifo0.fifo_store[81][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16109_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01248_),
    .Q(\fifo0.fifo_store[81][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16110_ (.CLK(clknet_leaf_210_clk_i),
    .D(_01249_),
    .Q(\fifo0.fifo_store[81][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16111_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01250_),
    .Q(\fifo0.fifo_store[81][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16112_ (.CLK(clknet_leaf_238_clk_i),
    .D(_01251_),
    .Q(\fifo0.fifo_store[81][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16113_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01252_),
    .Q(\fifo0.fifo_store[81][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16114_ (.CLK(clknet_leaf_238_clk_i),
    .D(_01253_),
    .Q(\fifo0.fifo_store[81][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16115_ (.CLK(clknet_leaf_215_clk_i),
    .D(_01254_),
    .Q(\fifo0.fifo_store[81][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16116_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01255_),
    .Q(\fifo0.fifo_store[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16117_ (.CLK(clknet_leaf_81_clk_i),
    .D(_01256_),
    .Q(\fifo0.fifo_store[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16118_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01257_),
    .Q(\fifo0.fifo_store[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16119_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01258_),
    .Q(\fifo0.fifo_store[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16120_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01259_),
    .Q(\fifo0.fifo_store[94][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16121_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01260_),
    .Q(\fifo0.fifo_store[94][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16122_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01261_),
    .Q(\fifo0.fifo_store[94][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16123_ (.CLK(clknet_leaf_151_clk_i),
    .D(_01262_),
    .Q(\fifo0.fifo_store[94][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16124_ (.CLK(clknet_leaf_135_clk_i),
    .D(_01263_),
    .Q(\fifo0.fifo_store[94][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16125_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01264_),
    .Q(\fifo0.fifo_store[94][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16126_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01265_),
    .Q(\fifo0.fifo_store[94][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16127_ (.CLK(clknet_leaf_176_clk_i),
    .D(_01266_),
    .Q(\fifo0.fifo_store[94][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16128_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01267_),
    .Q(\fifo0.fifo_store[94][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16129_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01268_),
    .Q(\fifo0.fifo_store[94][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16130_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01269_),
    .Q(\fifo0.fifo_store[94][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16131_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01270_),
    .Q(\fifo0.fifo_store[94][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16132_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01271_),
    .Q(\fifo0.fifo_store[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16133_ (.CLK(clknet_leaf_12_clk_i),
    .D(_01272_),
    .Q(\fifo0.fifo_store[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16134_ (.CLK(clknet_leaf_37_clk_i),
    .D(_01273_),
    .Q(\fifo0.fifo_store[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16135_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01274_),
    .Q(\fifo0.fifo_store[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16136_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01275_),
    .Q(\fifo0.fifo_store[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16137_ (.CLK(clknet_leaf_32_clk_i),
    .D(_01276_),
    .Q(\fifo0.fifo_store[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16138_ (.CLK(clknet_leaf_35_clk_i),
    .D(_01277_),
    .Q(\fifo0.fifo_store[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16139_ (.CLK(clknet_leaf_214_clk_i),
    .D(_01278_),
    .Q(\fifo0.fifo_store[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16140_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01279_),
    .Q(\fifo0.fifo_store[44][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16141_ (.CLK(clknet_leaf_39_clk_i),
    .D(_01280_),
    .Q(\fifo0.fifo_store[44][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16142_ (.CLK(clknet_leaf_229_clk_i),
    .D(_01281_),
    .Q(\fifo0.fifo_store[44][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16143_ (.CLK(clknet_leaf_249_clk_i),
    .D(_01282_),
    .Q(\fifo0.fifo_store[44][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16144_ (.CLK(clknet_leaf_240_clk_i),
    .D(_01283_),
    .Q(\fifo0.fifo_store[44][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16145_ (.CLK(clknet_leaf_244_clk_i),
    .D(_01284_),
    .Q(\fifo0.fifo_store[44][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16146_ (.CLK(clknet_leaf_239_clk_i),
    .D(_01285_),
    .Q(\fifo0.fifo_store[44][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16147_ (.CLK(clknet_leaf_292_clk_i),
    .D(_01286_),
    .Q(\fifo0.fifo_store[44][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16148_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01287_),
    .Q(\fifo0.fifo_store[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16149_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01288_),
    .Q(\fifo0.fifo_store[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16150_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01289_),
    .Q(\fifo0.fifo_store[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16151_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01290_),
    .Q(\fifo0.fifo_store[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16152_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01291_),
    .Q(\fifo0.fifo_store[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16153_ (.CLK(clknet_leaf_304_clk_i),
    .D(_01292_),
    .Q(\fifo0.fifo_store[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16154_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01293_),
    .Q(\fifo0.fifo_store[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16155_ (.CLK(clknet_leaf_299_clk_i),
    .D(_01294_),
    .Q(\fifo0.fifo_store[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16156_ (.CLK(clknet_leaf_306_clk_i),
    .D(_01295_),
    .Q(\fifo0.fifo_store[43][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16157_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01296_),
    .Q(\fifo0.fifo_store[43][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16158_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01297_),
    .Q(\fifo0.fifo_store[43][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16159_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01298_),
    .Q(\fifo0.fifo_store[43][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16160_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01299_),
    .Q(\fifo0.fifo_store[43][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16161_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01300_),
    .Q(\fifo0.fifo_store[43][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16162_ (.CLK(clknet_leaf_264_clk_i),
    .D(_01301_),
    .Q(\fifo0.fifo_store[43][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16163_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01302_),
    .Q(\fifo0.fifo_store[43][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16164_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01303_),
    .Q(\fifo0.fifo_store[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16165_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01304_),
    .Q(\fifo0.fifo_store[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16166_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01305_),
    .Q(\fifo0.fifo_store[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16167_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01306_),
    .Q(\fifo0.fifo_store[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16168_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01307_),
    .Q(\fifo0.fifo_store[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16169_ (.CLK(clknet_leaf_304_clk_i),
    .D(_01308_),
    .Q(\fifo0.fifo_store[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16170_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01309_),
    .Q(\fifo0.fifo_store[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16171_ (.CLK(clknet_leaf_298_clk_i),
    .D(_01310_),
    .Q(\fifo0.fifo_store[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16172_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01311_),
    .Q(\fifo0.fifo_store[42][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16173_ (.CLK(clknet_leaf_314_clk_i),
    .D(_01312_),
    .Q(\fifo0.fifo_store[42][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16174_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01313_),
    .Q(\fifo0.fifo_store[42][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16175_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01314_),
    .Q(\fifo0.fifo_store[42][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16176_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01315_),
    .Q(\fifo0.fifo_store[42][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16177_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01316_),
    .Q(\fifo0.fifo_store[42][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16178_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01317_),
    .Q(\fifo0.fifo_store[42][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16179_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01318_),
    .Q(\fifo0.fifo_store[42][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16180_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01319_),
    .Q(\fifo0.fifo_store[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16181_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01320_),
    .Q(\fifo0.fifo_store[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16182_ (.CLK(clknet_leaf_309_clk_i),
    .D(_01321_),
    .Q(\fifo0.fifo_store[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16183_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01322_),
    .Q(\fifo0.fifo_store[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16184_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01323_),
    .Q(\fifo0.fifo_store[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16185_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01324_),
    .Q(\fifo0.fifo_store[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16186_ (.CLK(clknet_leaf_310_clk_i),
    .D(_01325_),
    .Q(\fifo0.fifo_store[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16187_ (.CLK(clknet_leaf_298_clk_i),
    .D(_01326_),
    .Q(\fifo0.fifo_store[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16188_ (.CLK(clknet_leaf_297_clk_i),
    .D(_01327_),
    .Q(\fifo0.fifo_store[41][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16189_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01328_),
    .Q(\fifo0.fifo_store[41][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16190_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01329_),
    .Q(\fifo0.fifo_store[41][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16191_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01330_),
    .Q(\fifo0.fifo_store[41][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16192_ (.CLK(clknet_leaf_251_clk_i),
    .D(_01331_),
    .Q(\fifo0.fifo_store[41][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16193_ (.CLK(clknet_leaf_251_clk_i),
    .D(_01332_),
    .Q(\fifo0.fifo_store[41][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16194_ (.CLK(clknet_leaf_253_clk_i),
    .D(_01333_),
    .Q(\fifo0.fifo_store[41][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16195_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01334_),
    .Q(\fifo0.fifo_store[41][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16196_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01335_),
    .Q(\fifo0.fifo_store[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16197_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01336_),
    .Q(\fifo0.fifo_store[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16198_ (.CLK(clknet_leaf_309_clk_i),
    .D(_01337_),
    .Q(\fifo0.fifo_store[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16199_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01338_),
    .Q(\fifo0.fifo_store[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16200_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01339_),
    .Q(\fifo0.fifo_store[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16201_ (.CLK(clknet_leaf_304_clk_i),
    .D(_01340_),
    .Q(\fifo0.fifo_store[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16202_ (.CLK(clknet_leaf_310_clk_i),
    .D(_01341_),
    .Q(\fifo0.fifo_store[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16203_ (.CLK(clknet_leaf_297_clk_i),
    .D(_01342_),
    .Q(\fifo0.fifo_store[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16204_ (.CLK(clknet_leaf_306_clk_i),
    .D(_01343_),
    .Q(\fifo0.fifo_store[40][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16205_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01344_),
    .Q(\fifo0.fifo_store[40][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16206_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01345_),
    .Q(\fifo0.fifo_store[40][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16207_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01346_),
    .Q(\fifo0.fifo_store[40][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16208_ (.CLK(clknet_leaf_251_clk_i),
    .D(_01347_),
    .Q(\fifo0.fifo_store[40][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16209_ (.CLK(clknet_leaf_251_clk_i),
    .D(_01348_),
    .Q(\fifo0.fifo_store[40][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16210_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01349_),
    .Q(\fifo0.fifo_store[40][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16211_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01350_),
    .Q(\fifo0.fifo_store[40][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16212_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01351_),
    .Q(\fifo0.fifo_store[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16213_ (.CLK(clknet_leaf_13_clk_i),
    .D(_01352_),
    .Q(\fifo0.fifo_store[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16214_ (.CLK(clknet_leaf_29_clk_i),
    .D(_01353_),
    .Q(\fifo0.fifo_store[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16215_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01354_),
    .Q(\fifo0.fifo_store[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16216_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01355_),
    .Q(\fifo0.fifo_store[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16217_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01356_),
    .Q(\fifo0.fifo_store[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16218_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01357_),
    .Q(\fifo0.fifo_store[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16219_ (.CLK(clknet_leaf_299_clk_i),
    .D(_01358_),
    .Q(\fifo0.fifo_store[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16220_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01359_),
    .Q(\fifo0.fifo_store[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16221_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01360_),
    .Q(\fifo0.fifo_store[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16222_ (.CLK(clknet_leaf_226_clk_i),
    .D(_01361_),
    .Q(\fifo0.fifo_store[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16223_ (.CLK(clknet_leaf_227_clk_i),
    .D(_01362_),
    .Q(\fifo0.fifo_store[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16224_ (.CLK(clknet_leaf_228_clk_i),
    .D(_01363_),
    .Q(\fifo0.fifo_store[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16225_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01364_),
    .Q(\fifo0.fifo_store[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16226_ (.CLK(clknet_leaf_229_clk_i),
    .D(_01365_),
    .Q(\fifo0.fifo_store[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16227_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01366_),
    .Q(\fifo0.fifo_store[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16228_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01367_),
    .Q(\fifo0.fifo_store[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16229_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01368_),
    .Q(\fifo0.fifo_store[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16230_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01369_),
    .Q(\fifo0.fifo_store[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16231_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01370_),
    .Q(\fifo0.fifo_store[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16232_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01371_),
    .Q(\fifo0.fifo_store[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16233_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01372_),
    .Q(\fifo0.fifo_store[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16234_ (.CLK(clknet_leaf_309_clk_i),
    .D(_01373_),
    .Q(\fifo0.fifo_store[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16235_ (.CLK(clknet_leaf_298_clk_i),
    .D(_01374_),
    .Q(\fifo0.fifo_store[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16236_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01375_),
    .Q(\fifo0.fifo_store[38][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16237_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01376_),
    .Q(\fifo0.fifo_store[38][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16238_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01377_),
    .Q(\fifo0.fifo_store[38][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16239_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01378_),
    .Q(\fifo0.fifo_store[38][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16240_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01379_),
    .Q(\fifo0.fifo_store[38][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16241_ (.CLK(clknet_leaf_246_clk_i),
    .D(_01380_),
    .Q(\fifo0.fifo_store[38][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16242_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01381_),
    .Q(\fifo0.fifo_store[38][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16243_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01382_),
    .Q(\fifo0.fifo_store[38][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16244_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01383_),
    .Q(\fifo0.fifo_store[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16245_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01384_),
    .Q(\fifo0.fifo_store[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16246_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01385_),
    .Q(\fifo0.fifo_store[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16247_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01386_),
    .Q(\fifo0.fifo_store[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16248_ (.CLK(clknet_leaf_314_clk_i),
    .D(_01387_),
    .Q(\fifo0.fifo_store[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16249_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01388_),
    .Q(\fifo0.fifo_store[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16250_ (.CLK(clknet_leaf_308_clk_i),
    .D(_01389_),
    .Q(\fifo0.fifo_store[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16251_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01390_),
    .Q(\fifo0.fifo_store[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16252_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01391_),
    .Q(\fifo0.fifo_store[37][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16253_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01392_),
    .Q(\fifo0.fifo_store[37][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16254_ (.CLK(clknet_leaf_290_clk_i),
    .D(_01393_),
    .Q(\fifo0.fifo_store[37][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16255_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01394_),
    .Q(\fifo0.fifo_store[37][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16256_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01395_),
    .Q(\fifo0.fifo_store[37][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16257_ (.CLK(clknet_leaf_245_clk_i),
    .D(_01396_),
    .Q(\fifo0.fifo_store[37][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16258_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01397_),
    .Q(\fifo0.fifo_store[37][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16259_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01398_),
    .Q(\fifo0.fifo_store[37][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16260_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01399_),
    .Q(\fifo0.fifo_store[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16261_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01400_),
    .Q(\fifo0.fifo_store[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16262_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01401_),
    .Q(\fifo0.fifo_store[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16263_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01402_),
    .Q(\fifo0.fifo_store[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16264_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01403_),
    .Q(\fifo0.fifo_store[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16265_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01404_),
    .Q(\fifo0.fifo_store[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16266_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01405_),
    .Q(\fifo0.fifo_store[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16267_ (.CLK(clknet_leaf_220_clk_i),
    .D(_01406_),
    .Q(\fifo0.fifo_store[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16268_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01407_),
    .Q(\fifo0.fifo_store[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16269_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01408_),
    .Q(\fifo0.fifo_store[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16270_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01409_),
    .Q(\fifo0.fifo_store[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16271_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01410_),
    .Q(\fifo0.fifo_store[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16272_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01411_),
    .Q(\fifo0.fifo_store[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16273_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01412_),
    .Q(\fifo0.fifo_store[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16274_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01413_),
    .Q(\fifo0.fifo_store[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16275_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01414_),
    .Q(\fifo0.fifo_store[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16276_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01415_),
    .Q(\fifo0.fifo_store[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16277_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01416_),
    .Q(\fifo0.fifo_store[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16278_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01417_),
    .Q(\fifo0.fifo_store[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16279_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01418_),
    .Q(\fifo0.fifo_store[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16280_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01419_),
    .Q(\fifo0.fifo_store[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16281_ (.CLK(clknet_leaf_306_clk_i),
    .D(_01420_),
    .Q(\fifo0.fifo_store[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16282_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01421_),
    .Q(\fifo0.fifo_store[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16283_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01422_),
    .Q(\fifo0.fifo_store[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16284_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01423_),
    .Q(\fifo0.fifo_store[36][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16285_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01424_),
    .Q(\fifo0.fifo_store[36][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16286_ (.CLK(clknet_leaf_290_clk_i),
    .D(_01425_),
    .Q(\fifo0.fifo_store[36][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16287_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01426_),
    .Q(\fifo0.fifo_store[36][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16288_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01427_),
    .Q(\fifo0.fifo_store[36][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16289_ (.CLK(clknet_leaf_245_clk_i),
    .D(_01428_),
    .Q(\fifo0.fifo_store[36][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16290_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01429_),
    .Q(\fifo0.fifo_store[36][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16291_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01430_),
    .Q(\fifo0.fifo_store[36][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16292_ (.CLK(clknet_leaf_3_clk_i),
    .D(_01431_),
    .Q(\fifo0.fifo_store[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16293_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01432_),
    .Q(\fifo0.fifo_store[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16294_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01433_),
    .Q(\fifo0.fifo_store[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16295_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01434_),
    .Q(\fifo0.fifo_store[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16296_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01435_),
    .Q(\fifo0.fifo_store[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16297_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01436_),
    .Q(\fifo0.fifo_store[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16298_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01437_),
    .Q(\fifo0.fifo_store[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16299_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01438_),
    .Q(\fifo0.fifo_store[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16300_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01439_),
    .Q(\fifo0.fifo_store[35][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16301_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01440_),
    .Q(\fifo0.fifo_store[35][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16302_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01441_),
    .Q(\fifo0.fifo_store[35][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16303_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01442_),
    .Q(\fifo0.fifo_store[35][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16304_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01443_),
    .Q(\fifo0.fifo_store[35][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16305_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01444_),
    .Q(\fifo0.fifo_store[35][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16306_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01445_),
    .Q(\fifo0.fifo_store[35][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16307_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01446_),
    .Q(\fifo0.fifo_store[35][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16308_ (.CLK(clknet_leaf_3_clk_i),
    .D(_01447_),
    .Q(\fifo0.fifo_store[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16309_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01448_),
    .Q(\fifo0.fifo_store[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16310_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01449_),
    .Q(\fifo0.fifo_store[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16311_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01450_),
    .Q(\fifo0.fifo_store[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16312_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01451_),
    .Q(\fifo0.fifo_store[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16313_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01452_),
    .Q(\fifo0.fifo_store[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16314_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01453_),
    .Q(\fifo0.fifo_store[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16315_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01454_),
    .Q(\fifo0.fifo_store[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16316_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01455_),
    .Q(\fifo0.fifo_store[34][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16317_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01456_),
    .Q(\fifo0.fifo_store[34][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16318_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01457_),
    .Q(\fifo0.fifo_store[34][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16319_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01458_),
    .Q(\fifo0.fifo_store[34][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16320_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01459_),
    .Q(\fifo0.fifo_store[34][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16321_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01460_),
    .Q(\fifo0.fifo_store[34][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16322_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01461_),
    .Q(\fifo0.fifo_store[34][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16323_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01462_),
    .Q(\fifo0.fifo_store[34][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16324_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01463_),
    .Q(\fifo0.fifo_store[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16325_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01464_),
    .Q(\fifo0.fifo_store[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16326_ (.CLK(clknet_leaf_31_clk_i),
    .D(_01465_),
    .Q(\fifo0.fifo_store[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16327_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01466_),
    .Q(\fifo0.fifo_store[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16328_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01467_),
    .Q(\fifo0.fifo_store[99][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16329_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01468_),
    .Q(\fifo0.fifo_store[99][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16330_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01469_),
    .Q(\fifo0.fifo_store[99][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16331_ (.CLK(clknet_leaf_215_clk_i),
    .D(_01470_),
    .Q(\fifo0.fifo_store[99][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16332_ (.CLK(clknet_leaf_216_clk_i),
    .D(_01471_),
    .Q(\fifo0.fifo_store[99][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16333_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01472_),
    .Q(\fifo0.fifo_store[99][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16334_ (.CLK(clknet_leaf_227_clk_i),
    .D(_01473_),
    .Q(\fifo0.fifo_store[99][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16335_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01474_),
    .Q(\fifo0.fifo_store[99][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16336_ (.CLK(clknet_leaf_241_clk_i),
    .D(_01475_),
    .Q(\fifo0.fifo_store[99][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16337_ (.CLK(clknet_leaf_246_clk_i),
    .D(_01476_),
    .Q(\fifo0.fifo_store[99][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16338_ (.CLK(clknet_leaf_242_clk_i),
    .D(_01477_),
    .Q(\fifo0.fifo_store[99][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16339_ (.CLK(clknet_leaf_291_clk_i),
    .D(_01478_),
    .Q(\fifo0.fifo_store[99][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16340_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01479_),
    .Q(\fifo0.fifo_store[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16341_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01480_),
    .Q(\fifo0.fifo_store[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16342_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01481_),
    .Q(\fifo0.fifo_store[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16343_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01482_),
    .Q(\fifo0.fifo_store[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16344_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01483_),
    .Q(\fifo0.fifo_store[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16345_ (.CLK(clknet_leaf_283_clk_i),
    .D(_01484_),
    .Q(\fifo0.fifo_store[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16346_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01485_),
    .Q(\fifo0.fifo_store[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16347_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01486_),
    .Q(\fifo0.fifo_store[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16348_ (.CLK(clknet_leaf_306_clk_i),
    .D(_01487_),
    .Q(\fifo0.fifo_store[33][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16349_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01488_),
    .Q(\fifo0.fifo_store[33][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16350_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01489_),
    .Q(\fifo0.fifo_store[33][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16351_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01490_),
    .Q(\fifo0.fifo_store[33][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16352_ (.CLK(clknet_leaf_265_clk_i),
    .D(_01491_),
    .Q(\fifo0.fifo_store[33][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16353_ (.CLK(clknet_leaf_264_clk_i),
    .D(_01492_),
    .Q(\fifo0.fifo_store[33][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16354_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01493_),
    .Q(\fifo0.fifo_store[33][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16355_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01494_),
    .Q(\fifo0.fifo_store[33][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16356_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01495_),
    .Q(\fifo0.fifo_store[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16357_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01496_),
    .Q(\fifo0.fifo_store[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16358_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01497_),
    .Q(\fifo0.fifo_store[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16359_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01498_),
    .Q(\fifo0.fifo_store[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16360_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01499_),
    .Q(\fifo0.fifo_store[89][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16361_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01500_),
    .Q(\fifo0.fifo_store[89][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16362_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01501_),
    .Q(\fifo0.fifo_store[89][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16363_ (.CLK(clknet_leaf_141_clk_i),
    .D(_01502_),
    .Q(\fifo0.fifo_store[89][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16364_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01503_),
    .Q(\fifo0.fifo_store[89][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16365_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01504_),
    .Q(\fifo0.fifo_store[89][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16366_ (.CLK(clknet_leaf_206_clk_i),
    .D(_01505_),
    .Q(\fifo0.fifo_store[89][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16367_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01506_),
    .Q(\fifo0.fifo_store[89][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16368_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01507_),
    .Q(\fifo0.fifo_store[89][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16369_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01508_),
    .Q(\fifo0.fifo_store[89][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16370_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01509_),
    .Q(\fifo0.fifo_store[89][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16371_ (.CLK(clknet_leaf_208_clk_i),
    .D(_01510_),
    .Q(\fifo0.fifo_store[89][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16372_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01511_),
    .Q(\fifo0.fifo_store[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16373_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01512_),
    .Q(\fifo0.fifo_store[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16374_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01513_),
    .Q(\fifo0.fifo_store[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16375_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01514_),
    .Q(\fifo0.fifo_store[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16376_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01515_),
    .Q(\fifo0.fifo_store[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16377_ (.CLK(clknet_leaf_283_clk_i),
    .D(_01516_),
    .Q(\fifo0.fifo_store[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16378_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01517_),
    .Q(\fifo0.fifo_store[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16379_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01518_),
    .Q(\fifo0.fifo_store[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16380_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01519_),
    .Q(\fifo0.fifo_store[32][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16381_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01520_),
    .Q(\fifo0.fifo_store[32][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16382_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01521_),
    .Q(\fifo0.fifo_store[32][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16383_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01522_),
    .Q(\fifo0.fifo_store[32][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16384_ (.CLK(clknet_leaf_264_clk_i),
    .D(_01523_),
    .Q(\fifo0.fifo_store[32][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16385_ (.CLK(clknet_leaf_264_clk_i),
    .D(_01524_),
    .Q(\fifo0.fifo_store[32][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16386_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01525_),
    .Q(\fifo0.fifo_store[32][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16387_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01526_),
    .Q(\fifo0.fifo_store[32][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16388_ (.CLK(clknet_leaf_3_clk_i),
    .D(_01527_),
    .Q(\fifo0.fifo_store[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16389_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01528_),
    .Q(\fifo0.fifo_store[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16390_ (.CLK(clknet_leaf_321_clk_i),
    .D(_01529_),
    .Q(\fifo0.fifo_store[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16391_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01530_),
    .Q(\fifo0.fifo_store[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16392_ (.CLK(clknet_leaf_333_clk_i),
    .D(_01531_),
    .Q(\fifo0.fifo_store[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16393_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01532_),
    .Q(\fifo0.fifo_store[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16394_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01533_),
    .Q(\fifo0.fifo_store[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16395_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01534_),
    .Q(\fifo0.fifo_store[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16396_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01535_),
    .Q(\fifo0.fifo_store[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16397_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01536_),
    .Q(\fifo0.fifo_store[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16398_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01537_),
    .Q(\fifo0.fifo_store[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16399_ (.CLK(clknet_leaf_267_clk_i),
    .D(_01538_),
    .Q(\fifo0.fifo_store[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16400_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01539_),
    .Q(\fifo0.fifo_store[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16401_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01540_),
    .Q(\fifo0.fifo_store[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16402_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01541_),
    .Q(\fifo0.fifo_store[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16403_ (.CLK(clknet_leaf_281_clk_i),
    .D(_01542_),
    .Q(\fifo0.fifo_store[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16404_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01543_),
    .Q(\fifo0.fifo_store[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16405_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01544_),
    .Q(\fifo0.fifo_store[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16406_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01545_),
    .Q(\fifo0.fifo_store[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16407_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01546_),
    .Q(\fifo0.fifo_store[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16408_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01547_),
    .Q(\fifo0.fifo_store[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16409_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01548_),
    .Q(\fifo0.fifo_store[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16410_ (.CLK(clknet_leaf_315_clk_i),
    .D(_01549_),
    .Q(\fifo0.fifo_store[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16411_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01550_),
    .Q(\fifo0.fifo_store[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16412_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01551_),
    .Q(\fifo0.fifo_store[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16413_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01552_),
    .Q(\fifo0.fifo_store[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16414_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01553_),
    .Q(\fifo0.fifo_store[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16415_ (.CLK(clknet_leaf_267_clk_i),
    .D(_01554_),
    .Q(\fifo0.fifo_store[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16416_ (.CLK(clknet_leaf_253_clk_i),
    .D(_01555_),
    .Q(\fifo0.fifo_store[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16417_ (.CLK(clknet_leaf_252_clk_i),
    .D(_01556_),
    .Q(\fifo0.fifo_store[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16418_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01557_),
    .Q(\fifo0.fifo_store[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16419_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01558_),
    .Q(\fifo0.fifo_store[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16420_ (.CLK(clknet_leaf_3_clk_i),
    .D(_01559_),
    .Q(\fifo0.fifo_store[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16421_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01560_),
    .Q(\fifo0.fifo_store[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16422_ (.CLK(clknet_leaf_321_clk_i),
    .D(_01561_),
    .Q(\fifo0.fifo_store[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16423_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01562_),
    .Q(\fifo0.fifo_store[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16424_ (.CLK(clknet_leaf_333_clk_i),
    .D(_01563_),
    .Q(\fifo0.fifo_store[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16425_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01564_),
    .Q(\fifo0.fifo_store[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16426_ (.CLK(clknet_leaf_317_clk_i),
    .D(_01565_),
    .Q(\fifo0.fifo_store[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16427_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01566_),
    .Q(\fifo0.fifo_store[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16428_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01567_),
    .Q(\fifo0.fifo_store[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16429_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01568_),
    .Q(\fifo0.fifo_store[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16430_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01569_),
    .Q(\fifo0.fifo_store[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16431_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01570_),
    .Q(\fifo0.fifo_store[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16432_ (.CLK(clknet_leaf_253_clk_i),
    .D(_01571_),
    .Q(\fifo0.fifo_store[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16433_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01572_),
    .Q(\fifo0.fifo_store[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16434_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01573_),
    .Q(\fifo0.fifo_store[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16435_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01574_),
    .Q(\fifo0.fifo_store[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16436_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01575_),
    .Q(\fifo0.fifo_store[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16437_ (.CLK(clknet_leaf_13_clk_i),
    .D(_01576_),
    .Q(\fifo0.fifo_store[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16438_ (.CLK(clknet_leaf_29_clk_i),
    .D(_01577_),
    .Q(\fifo0.fifo_store[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16439_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01578_),
    .Q(\fifo0.fifo_store[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16440_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01579_),
    .Q(\fifo0.fifo_store[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16441_ (.CLK(clknet_leaf_301_clk_i),
    .D(_01580_),
    .Q(\fifo0.fifo_store[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16442_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01581_),
    .Q(\fifo0.fifo_store[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16443_ (.CLK(clknet_leaf_299_clk_i),
    .D(_01582_),
    .Q(\fifo0.fifo_store[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16444_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01583_),
    .Q(\fifo0.fifo_store[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16445_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01584_),
    .Q(\fifo0.fifo_store[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16446_ (.CLK(clknet_leaf_226_clk_i),
    .D(_01585_),
    .Q(\fifo0.fifo_store[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16447_ (.CLK(clknet_leaf_227_clk_i),
    .D(_01586_),
    .Q(\fifo0.fifo_store[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16448_ (.CLK(clknet_leaf_228_clk_i),
    .D(_01587_),
    .Q(\fifo0.fifo_store[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16449_ (.CLK(clknet_leaf_250_clk_i),
    .D(_01588_),
    .Q(\fifo0.fifo_store[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16450_ (.CLK(clknet_leaf_229_clk_i),
    .D(_01589_),
    .Q(\fifo0.fifo_store[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16451_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01590_),
    .Q(\fifo0.fifo_store[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16452_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01591_),
    .Q(\fifo0.fifo_store[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16453_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01592_),
    .Q(\fifo0.fifo_store[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16454_ (.CLK(clknet_leaf_317_clk_i),
    .D(_01593_),
    .Q(\fifo0.fifo_store[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16455_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01594_),
    .Q(\fifo0.fifo_store[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16456_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01595_),
    .Q(\fifo0.fifo_store[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16457_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01596_),
    .Q(\fifo0.fifo_store[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16458_ (.CLK(clknet_leaf_311_clk_i),
    .D(_01597_),
    .Q(\fifo0.fifo_store[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16459_ (.CLK(clknet_leaf_299_clk_i),
    .D(_01598_),
    .Q(\fifo0.fifo_store[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16460_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01599_),
    .Q(\fifo0.fifo_store[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16461_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01600_),
    .Q(\fifo0.fifo_store[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16462_ (.CLK(clknet_leaf_267_clk_i),
    .D(_01601_),
    .Q(\fifo0.fifo_store[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16463_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01602_),
    .Q(\fifo0.fifo_store[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16464_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01603_),
    .Q(\fifo0.fifo_store[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16465_ (.CLK(clknet_leaf_244_clk_i),
    .D(_01604_),
    .Q(\fifo0.fifo_store[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16466_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01605_),
    .Q(\fifo0.fifo_store[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16467_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01606_),
    .Q(\fifo0.fifo_store[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16468_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01607_),
    .Q(\fifo0.fifo_store[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16469_ (.CLK(clknet_leaf_15_clk_i),
    .D(_01608_),
    .Q(\fifo0.fifo_store[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16470_ (.CLK(clknet_leaf_304_clk_i),
    .D(_01609_),
    .Q(\fifo0.fifo_store[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16471_ (.CLK(clknet_leaf_16_clk_i),
    .D(_01610_),
    .Q(\fifo0.fifo_store[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16472_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01611_),
    .Q(\fifo0.fifo_store[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16473_ (.CLK(clknet_leaf_301_clk_i),
    .D(_01612_),
    .Q(\fifo0.fifo_store[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16474_ (.CLK(clknet_leaf_30_clk_i),
    .D(_01613_),
    .Q(\fifo0.fifo_store[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16475_ (.CLK(clknet_leaf_220_clk_i),
    .D(_01614_),
    .Q(\fifo0.fifo_store[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16476_ (.CLK(clknet_leaf_302_clk_i),
    .D(_01615_),
    .Q(\fifo0.fifo_store[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16477_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01616_),
    .Q(\fifo0.fifo_store[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16478_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01617_),
    .Q(\fifo0.fifo_store[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16479_ (.CLK(clknet_leaf_232_clk_i),
    .D(_01618_),
    .Q(\fifo0.fifo_store[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16480_ (.CLK(clknet_leaf_231_clk_i),
    .D(_01619_),
    .Q(\fifo0.fifo_store[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16481_ (.CLK(clknet_leaf_231_clk_i),
    .D(_01620_),
    .Q(\fifo0.fifo_store[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16482_ (.CLK(clknet_leaf_230_clk_i),
    .D(_01621_),
    .Q(\fifo0.fifo_store[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16483_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01622_),
    .Q(\fifo0.fifo_store[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16484_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01623_),
    .Q(\fifo0.fifo_data_del1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16485_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01624_),
    .Q(\fifo0.fifo_data_del1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16486_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01625_),
    .Q(\fifo0.fifo_data_del1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16487_ (.CLK(clknet_leaf_337_clk_i),
    .D(_01626_),
    .Q(\fifo0.fifo_data_del1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16488_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01627_),
    .Q(\fifo0.fifo_data_del1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16489_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01628_),
    .Q(\fifo0.fifo_data_del1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _16490_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01629_),
    .Q(\fifo0.fifo_data_del1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16491_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01630_),
    .Q(\fifo0.fifo_data_del1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _16492_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01631_),
    .Q(\fifo0.fifo_data_del1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _16493_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01632_),
    .Q(\fifo0.fifo_data_del1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _16494_ (.CLK(clknet_leaf_278_clk_i),
    .D(_01633_),
    .Q(\fifo0.fifo_data_del1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _16495_ (.CLK(clknet_leaf_278_clk_i),
    .D(_01634_),
    .Q(\fifo0.fifo_data_del1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _16496_ (.CLK(clknet_leaf_278_clk_i),
    .D(_01635_),
    .Q(\fifo0.fifo_data_del1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _16497_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01636_),
    .Q(\fifo0.fifo_data_del1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _16498_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01637_),
    .Q(\fifo0.fifo_data_del1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _16499_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01638_),
    .Q(\fifo0.fifo_data_del1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _16500_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01639_),
    .Q(\fifo0.fifo_rdy ));
 sky130_fd_sc_hd__dfxtp_1 _16501_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01640_),
    .Q(\fifo0.fifo_rdy_del1 ));
 sky130_fd_sc_hd__dfxtp_1 _16502_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01641_),
    .Q(\dsmod0.fetch_ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16503_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01642_),
    .Q(\dsmod0.fetch_ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16504_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01643_),
    .Q(\dsmod0.fetch_ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16505_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01644_),
    .Q(\dsmod0.fetch_ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16506_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01645_),
    .Q(\dsmod0.fetch_ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16507_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01646_),
    .Q(\dsmod0.fetch_ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _16508_ (.CLK(clknet_leaf_339_clk_i),
    .D(_01647_),
    .Q(\dsmod0.fetch_ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16509_ (.CLK(clknet_leaf_340_clk_i),
    .D(_01648_),
    .Q(\dsmod0.fetch_ctr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _16510_ (.CLK(clknet_5_16_0_clk_i),
    .D(_01649_),
    .Q(\fifo0.write_ptr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16511_ (.CLK(clknet_leaf_273_clk_i),
    .D(_01650_),
    .Q(\fifo0.write_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16512_ (.CLK(clknet_leaf_273_clk_i),
    .D(_01651_),
    .Q(\fifo0.write_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16513_ (.CLK(clknet_leaf_275_clk_i),
    .D(_01652_),
    .Q(\fifo0.write_ptr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16514_ (.CLK(clknet_leaf_275_clk_i),
    .D(_01653_),
    .Q(\fifo0.write_ptr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16515_ (.CLK(clknet_leaf_273_clk_i),
    .D(_01654_),
    .Q(\fifo0.write_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _16516_ (.CLK(clknet_leaf_277_clk_i),
    .D(_01655_),
    .Q(\fifo0.write_ptr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16517_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01656_),
    .Q(\fifo0.read_ptr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16518_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01657_),
    .Q(\fifo0.read_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16519_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01658_),
    .Q(\fifo0.read_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16520_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01659_),
    .Q(\fifo0.read_ptr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16521_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01660_),
    .Q(\fifo0.read_ptr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16522_ (.CLK(clknet_leaf_277_clk_i),
    .D(_01661_),
    .Q(\fifo0.read_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _16523_ (.CLK(clknet_leaf_277_clk_i),
    .D(_01662_),
    .Q(\fifo0.read_ptr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16524_ (.CLK(clknet_leaf_273_clk_i),
    .D(_01663_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _16525_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01664_),
    .Q(\fifo0.fifo_store[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16526_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01665_),
    .Q(\fifo0.fifo_store[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16527_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01666_),
    .Q(\fifo0.fifo_store[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16528_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01667_),
    .Q(\fifo0.fifo_store[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16529_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01668_),
    .Q(\fifo0.fifo_store[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16530_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01669_),
    .Q(\fifo0.fifo_store[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16531_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01670_),
    .Q(\fifo0.fifo_store[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16532_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01671_),
    .Q(\fifo0.fifo_store[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16533_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01672_),
    .Q(\fifo0.fifo_store[59][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16534_ (.CLK(clknet_leaf_39_clk_i),
    .D(_01673_),
    .Q(\fifo0.fifo_store[59][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16535_ (.CLK(clknet_leaf_223_clk_i),
    .D(_01674_),
    .Q(\fifo0.fifo_store[59][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16536_ (.CLK(clknet_leaf_234_clk_i),
    .D(_01675_),
    .Q(\fifo0.fifo_store[59][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16537_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01676_),
    .Q(\fifo0.fifo_store[59][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16538_ (.CLK(clknet_leaf_236_clk_i),
    .D(_01677_),
    .Q(\fifo0.fifo_store[59][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16539_ (.CLK(clknet_leaf_237_clk_i),
    .D(_01678_),
    .Q(\fifo0.fifo_store[59][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16540_ (.CLK(clknet_leaf_220_clk_i),
    .D(_01679_),
    .Q(\fifo0.fifo_store[59][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16541_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01680_),
    .Q(\fifo0.fifo_store[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16542_ (.CLK(clknet_leaf_13_clk_i),
    .D(_01681_),
    .Q(\fifo0.fifo_store[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16543_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01682_),
    .Q(\fifo0.fifo_store[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16544_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01683_),
    .Q(\fifo0.fifo_store[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16545_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01684_),
    .Q(\fifo0.fifo_store[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16546_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01685_),
    .Q(\fifo0.fifo_store[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16547_ (.CLK(clknet_leaf_310_clk_i),
    .D(_01686_),
    .Q(\fifo0.fifo_store[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16548_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01687_),
    .Q(\fifo0.fifo_store[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16549_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01688_),
    .Q(\fifo0.fifo_store[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16550_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01689_),
    .Q(\fifo0.fifo_store[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16551_ (.CLK(clknet_leaf_266_clk_i),
    .D(_01690_),
    .Q(\fifo0.fifo_store[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16552_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01691_),
    .Q(\fifo0.fifo_store[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16553_ (.CLK(clknet_leaf_255_clk_i),
    .D(_01692_),
    .Q(\fifo0.fifo_store[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16554_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01693_),
    .Q(\fifo0.fifo_store[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16555_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01694_),
    .Q(\fifo0.fifo_store[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16556_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01695_),
    .Q(\fifo0.fifo_store[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16557_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01696_),
    .Q(\fifo0.fifo_store[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16558_ (.CLK(clknet_leaf_4_clk_i),
    .D(_01697_),
    .Q(\fifo0.fifo_store[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16559_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01698_),
    .Q(\fifo0.fifo_store[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16560_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01699_),
    .Q(\fifo0.fifo_store[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16561_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01700_),
    .Q(\fifo0.fifo_store[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16562_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01701_),
    .Q(\fifo0.fifo_store[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16563_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01702_),
    .Q(\fifo0.fifo_store[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16564_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01703_),
    .Q(\fifo0.fifo_store[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16565_ (.CLK(clknet_leaf_308_clk_i),
    .D(_01704_),
    .Q(\fifo0.fifo_store[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16566_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01705_),
    .Q(\fifo0.fifo_store[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16567_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01706_),
    .Q(\fifo0.fifo_store[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16568_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01707_),
    .Q(\fifo0.fifo_store[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16569_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01708_),
    .Q(\fifo0.fifo_store[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16570_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01709_),
    .Q(\fifo0.fifo_store[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16571_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01710_),
    .Q(\fifo0.fifo_store[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16572_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01711_),
    .Q(\fifo0.fifo_store[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16573_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01712_),
    .Q(\fifo0.fifo_store[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16574_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01713_),
    .Q(\fifo0.fifo_store[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16575_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01714_),
    .Q(\fifo0.fifo_store[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16576_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01715_),
    .Q(\fifo0.fifo_store[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16577_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01716_),
    .Q(\fifo0.fifo_store[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16578_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01717_),
    .Q(\fifo0.fifo_store[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16579_ (.CLK(clknet_leaf_331_clk_i),
    .D(_01718_),
    .Q(\fifo0.fifo_store[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16580_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01719_),
    .Q(\fifo0.fifo_store[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16581_ (.CLK(clknet_leaf_308_clk_i),
    .D(_01720_),
    .Q(\fifo0.fifo_store[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16582_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01721_),
    .Q(\fifo0.fifo_store[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16583_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01722_),
    .Q(\fifo0.fifo_store[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16584_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01723_),
    .Q(\fifo0.fifo_store[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16585_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01724_),
    .Q(\fifo0.fifo_store[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16586_ (.CLK(clknet_leaf_260_clk_i),
    .D(_01725_),
    .Q(\fifo0.fifo_store[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16587_ (.CLK(clknet_leaf_260_clk_i),
    .D(_01726_),
    .Q(\fifo0.fifo_store[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16588_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01727_),
    .Q(\fifo0.fifo_store[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16589_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01728_),
    .Q(\fifo0.fifo_store[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16590_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01729_),
    .Q(\fifo0.fifo_store[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16591_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01730_),
    .Q(\fifo0.fifo_store[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16592_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01731_),
    .Q(\fifo0.fifo_store[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16593_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01732_),
    .Q(\fifo0.fifo_store[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16594_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01733_),
    .Q(\fifo0.fifo_store[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16595_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01734_),
    .Q(\fifo0.fifo_store[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16596_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01735_),
    .Q(\fifo0.fifo_store[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16597_ (.CLK(clknet_leaf_33_clk_i),
    .D(_01736_),
    .Q(\fifo0.fifo_store[48][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16598_ (.CLK(clknet_leaf_39_clk_i),
    .D(_01737_),
    .Q(\fifo0.fifo_store[48][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16599_ (.CLK(clknet_leaf_223_clk_i),
    .D(_01738_),
    .Q(\fifo0.fifo_store[48][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16600_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01739_),
    .Q(\fifo0.fifo_store[48][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16601_ (.CLK(clknet_leaf_235_clk_i),
    .D(_01740_),
    .Q(\fifo0.fifo_store[48][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16602_ (.CLK(clknet_leaf_234_clk_i),
    .D(_01741_),
    .Q(\fifo0.fifo_store[48][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16603_ (.CLK(clknet_leaf_233_clk_i),
    .D(_01742_),
    .Q(\fifo0.fifo_store[48][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16604_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01743_),
    .Q(\fifo0.fifo_store[48][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16605_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01744_),
    .Q(\fifo0.fifo_store[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16606_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01745_),
    .Q(\fifo0.fifo_store[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16607_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01746_),
    .Q(\fifo0.fifo_store[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16608_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01747_),
    .Q(\fifo0.fifo_store[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16609_ (.CLK(clknet_leaf_333_clk_i),
    .D(_01748_),
    .Q(\fifo0.fifo_store[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16610_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01749_),
    .Q(\fifo0.fifo_store[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16611_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01750_),
    .Q(\fifo0.fifo_store[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16612_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01751_),
    .Q(\fifo0.fifo_store[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16613_ (.CLK(clknet_leaf_309_clk_i),
    .D(_01752_),
    .Q(\fifo0.fifo_store[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16614_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01753_),
    .Q(\fifo0.fifo_store[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16615_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01754_),
    .Q(\fifo0.fifo_store[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16616_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01755_),
    .Q(\fifo0.fifo_store[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16617_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01756_),
    .Q(\fifo0.fifo_store[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16618_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01757_),
    .Q(\fifo0.fifo_store[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16619_ (.CLK(clknet_leaf_260_clk_i),
    .D(_01758_),
    .Q(\fifo0.fifo_store[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16620_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01759_),
    .Q(\fifo0.fifo_store[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16621_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01760_),
    .Q(\fifo0.fifo_store[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16622_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01761_),
    .Q(\fifo0.fifo_store[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16623_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01762_),
    .Q(\fifo0.fifo_store[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16624_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01763_),
    .Q(\fifo0.fifo_store[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16625_ (.CLK(clknet_leaf_314_clk_i),
    .D(_01764_),
    .Q(\fifo0.fifo_store[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16626_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01765_),
    .Q(\fifo0.fifo_store[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16627_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01766_),
    .Q(\fifo0.fifo_store[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16628_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01767_),
    .Q(\fifo0.fifo_store[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16629_ (.CLK(clknet_leaf_308_clk_i),
    .D(_01768_),
    .Q(\fifo0.fifo_store[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16630_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01769_),
    .Q(\fifo0.fifo_store[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16631_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01770_),
    .Q(\fifo0.fifo_store[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16632_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01771_),
    .Q(\fifo0.fifo_store[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16633_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01772_),
    .Q(\fifo0.fifo_store[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16634_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01773_),
    .Q(\fifo0.fifo_store[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16635_ (.CLK(clknet_leaf_260_clk_i),
    .D(_01774_),
    .Q(\fifo0.fifo_store[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16636_ (.CLK(clknet_leaf_269_clk_i),
    .D(_01775_),
    .Q(\fifo0.fifo_store[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16637_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01776_),
    .Q(\fifo0.fifo_store[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16638_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01777_),
    .Q(\fifo0.fifo_store[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16639_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01778_),
    .Q(\fifo0.fifo_store[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16640_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01779_),
    .Q(\fifo0.fifo_store[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16641_ (.CLK(clknet_leaf_314_clk_i),
    .D(_01780_),
    .Q(\fifo0.fifo_store[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16642_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01781_),
    .Q(\fifo0.fifo_store[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16643_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01782_),
    .Q(\fifo0.fifo_store[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16644_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01783_),
    .Q(\fifo0.fifo_store[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16645_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01784_),
    .Q(\fifo0.fifo_store[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16646_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01785_),
    .Q(\fifo0.fifo_store[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16647_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01786_),
    .Q(\fifo0.fifo_store[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16648_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01787_),
    .Q(\fifo0.fifo_store[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16649_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01788_),
    .Q(\fifo0.fifo_store[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16650_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01789_),
    .Q(\fifo0.fifo_store[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16651_ (.CLK(clknet_leaf_260_clk_i),
    .D(_01790_),
    .Q(\fifo0.fifo_store[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16652_ (.CLK(clknet_leaf_269_clk_i),
    .D(_01791_),
    .Q(\fifo0.fifo_store[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16653_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01792_),
    .Q(\fifo0.fifo_store[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16654_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01793_),
    .Q(\fifo0.fifo_store[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16655_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01794_),
    .Q(\fifo0.fifo_store[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16656_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01795_),
    .Q(\fifo0.fifo_store[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16657_ (.CLK(clknet_leaf_314_clk_i),
    .D(_01796_),
    .Q(\fifo0.fifo_store[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16658_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01797_),
    .Q(\fifo0.fifo_store[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16659_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01798_),
    .Q(\fifo0.fifo_store[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16660_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01799_),
    .Q(\fifo0.fifo_store[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16661_ (.CLK(clknet_leaf_310_clk_i),
    .D(_01800_),
    .Q(\fifo0.fifo_store[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16662_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01801_),
    .Q(\fifo0.fifo_store[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16663_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01802_),
    .Q(\fifo0.fifo_store[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16664_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01803_),
    .Q(\fifo0.fifo_store[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16665_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01804_),
    .Q(\fifo0.fifo_store[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16666_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01805_),
    .Q(\fifo0.fifo_store[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16667_ (.CLK(clknet_leaf_259_clk_i),
    .D(_01806_),
    .Q(\fifo0.fifo_store[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16668_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01807_),
    .Q(\fifo0.fifo_store[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16669_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01808_),
    .Q(\fifo0.fifo_store[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16670_ (.CLK(clknet_leaf_9_clk_i),
    .D(_01809_),
    .Q(\fifo0.fifo_store[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16671_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01810_),
    .Q(\fifo0.fifo_store[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16672_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01811_),
    .Q(\fifo0.fifo_store[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16673_ (.CLK(clknet_leaf_331_clk_i),
    .D(_01812_),
    .Q(\fifo0.fifo_store[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16674_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01813_),
    .Q(\fifo0.fifo_store[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16675_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01814_),
    .Q(\fifo0.fifo_store[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16676_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01815_),
    .Q(\fifo0.fifo_store[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16677_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01816_),
    .Q(\fifo0.fifo_store[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16678_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01817_),
    .Q(\fifo0.fifo_store[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16679_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01818_),
    .Q(\fifo0.fifo_store[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16680_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01819_),
    .Q(\fifo0.fifo_store[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16681_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01820_),
    .Q(\fifo0.fifo_store[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16682_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01821_),
    .Q(\fifo0.fifo_store[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16683_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01822_),
    .Q(\fifo0.fifo_store[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16684_ (.CLK(clknet_leaf_269_clk_i),
    .D(_01823_),
    .Q(\fifo0.fifo_store[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16685_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01824_),
    .Q(\fifo0.fifo_store[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16686_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01825_),
    .Q(\fifo0.fifo_store[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16687_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01826_),
    .Q(\fifo0.fifo_store[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16688_ (.CLK(clknet_leaf_342_clk_i),
    .D(_01827_),
    .Q(\fifo0.fifo_store[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16689_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01828_),
    .Q(\fifo0.fifo_store[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16690_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01829_),
    .Q(\fifo0.fifo_store[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16691_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01830_),
    .Q(\fifo0.fifo_store[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16692_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01831_),
    .Q(\fifo0.fifo_store[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16693_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01832_),
    .Q(\fifo0.fifo_store[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16694_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01833_),
    .Q(\fifo0.fifo_store[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16695_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01834_),
    .Q(\fifo0.fifo_store[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16696_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01835_),
    .Q(\fifo0.fifo_store[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16697_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01836_),
    .Q(\fifo0.fifo_store[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16698_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01837_),
    .Q(\fifo0.fifo_store[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16699_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01838_),
    .Q(\fifo0.fifo_store[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16700_ (.CLK(clknet_leaf_269_clk_i),
    .D(_01839_),
    .Q(\fifo0.fifo_store[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16701_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01840_),
    .Q(\fifo0.fifo_store[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16702_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01841_),
    .Q(\fifo0.fifo_store[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16703_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01842_),
    .Q(\fifo0.fifo_store[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16704_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01843_),
    .Q(\fifo0.fifo_store[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16705_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01844_),
    .Q(\fifo0.fifo_store[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16706_ (.CLK(clknet_leaf_297_clk_i),
    .D(_01845_),
    .Q(\fifo0.fifo_store[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16707_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01846_),
    .Q(\fifo0.fifo_store[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16708_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01847_),
    .Q(\fifo0.fifo_store[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16709_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01848_),
    .Q(\fifo0.fifo_store[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16710_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01849_),
    .Q(\fifo0.fifo_store[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16711_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01850_),
    .Q(\fifo0.fifo_store[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16712_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01851_),
    .Q(\fifo0.fifo_store[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16713_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01852_),
    .Q(\fifo0.fifo_store[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16714_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01853_),
    .Q(\fifo0.fifo_store[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16715_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01854_),
    .Q(\fifo0.fifo_store[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16716_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01855_),
    .Q(\fifo0.fifo_store[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16717_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01856_),
    .Q(\fifo0.fifo_store[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16718_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01857_),
    .Q(\fifo0.fifo_store[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16719_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01858_),
    .Q(\fifo0.fifo_store[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16720_ (.CLK(clknet_leaf_343_clk_i),
    .D(_01859_),
    .Q(\fifo0.fifo_store[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16721_ (.CLK(clknet_leaf_331_clk_i),
    .D(_01860_),
    .Q(\fifo0.fifo_store[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16722_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01861_),
    .Q(\fifo0.fifo_store[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16723_ (.CLK(clknet_leaf_321_clk_i),
    .D(_01862_),
    .Q(\fifo0.fifo_store[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16724_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01863_),
    .Q(\fifo0.fifo_store[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16725_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01864_),
    .Q(\fifo0.fifo_store[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16726_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01865_),
    .Q(\fifo0.fifo_store[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16727_ (.CLK(clknet_leaf_268_clk_i),
    .D(_01866_),
    .Q(\fifo0.fifo_store[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16728_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01867_),
    .Q(\fifo0.fifo_store[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16729_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01868_),
    .Q(\fifo0.fifo_store[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16730_ (.CLK(clknet_leaf_257_clk_i),
    .D(_01869_),
    .Q(\fifo0.fifo_store[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16731_ (.CLK(clknet_leaf_258_clk_i),
    .D(_01870_),
    .Q(\fifo0.fifo_store[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16732_ (.CLK(clknet_leaf_269_clk_i),
    .D(_01871_),
    .Q(\fifo0.fifo_store[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16733_ (.CLK(clknet_leaf_13_clk_i),
    .D(_01872_),
    .Q(\fifo0.fifo_store[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16734_ (.CLK(clknet_leaf_13_clk_i),
    .D(_01873_),
    .Q(\fifo0.fifo_store[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16735_ (.CLK(clknet_leaf_304_clk_i),
    .D(_01874_),
    .Q(\fifo0.fifo_store[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16736_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01875_),
    .Q(\fifo0.fifo_store[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16737_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01876_),
    .Q(\fifo0.fifo_store[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16738_ (.CLK(clknet_leaf_301_clk_i),
    .D(_01877_),
    .Q(\fifo0.fifo_store[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16739_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01878_),
    .Q(\fifo0.fifo_store[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16740_ (.CLK(clknet_leaf_219_clk_i),
    .D(_01879_),
    .Q(\fifo0.fifo_store[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16741_ (.CLK(clknet_leaf_303_clk_i),
    .D(_01880_),
    .Q(\fifo0.fifo_store[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16742_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01881_),
    .Q(\fifo0.fifo_store[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16743_ (.CLK(clknet_leaf_226_clk_i),
    .D(_01882_),
    .Q(\fifo0.fifo_store[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16744_ (.CLK(clknet_leaf_227_clk_i),
    .D(_01883_),
    .Q(\fifo0.fifo_store[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16745_ (.CLK(clknet_leaf_248_clk_i),
    .D(_01884_),
    .Q(\fifo0.fifo_store[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16746_ (.CLK(clknet_leaf_249_clk_i),
    .D(_01885_),
    .Q(\fifo0.fifo_store[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16747_ (.CLK(clknet_leaf_229_clk_i),
    .D(_01886_),
    .Q(\fifo0.fifo_store[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16748_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01887_),
    .Q(\fifo0.fifo_store[1][15] ));
 sky130_fd_sc_hd__dfxtp_4 _16749_ (.CLK(clknet_leaf_337_clk_i),
    .D(_01888_),
    .Q(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__dfxtp_4 _16750_ (.CLK(clknet_leaf_337_clk_i),
    .D(_01889_),
    .Q(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__dfxtp_4 _16751_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01890_),
    .Q(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__dfxtp_4 _16752_ (.CLK(clknet_leaf_337_clk_i),
    .D(_01891_),
    .Q(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__dfxtp_4 _16753_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01892_),
    .Q(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16754_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01893_),
    .Q(\fifo0.fifo_data[5] ));
 sky130_fd_sc_hd__dfxtp_4 _16755_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01894_),
    .Q(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16756_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01895_),
    .Q(\fifo0.fifo_data[7] ));
 sky130_fd_sc_hd__dfxtp_4 _16757_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01896_),
    .Q(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__dfxtp_4 _16758_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01897_),
    .Q(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _16759_ (.CLK(clknet_leaf_278_clk_i),
    .D(_01898_),
    .Q(\fifo0.fifo_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _16760_ (.CLK(clknet_leaf_278_clk_i),
    .D(_01899_),
    .Q(\fifo0.fifo_data[11] ));
 sky130_fd_sc_hd__dfxtp_4 _16761_ (.CLK(clknet_leaf_280_clk_i),
    .D(_01900_),
    .Q(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__dfxtp_4 _16762_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01901_),
    .Q(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__dfxtp_4 _16763_ (.CLK(clknet_leaf_271_clk_i),
    .D(_01902_),
    .Q(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__dfxtp_4 _16764_ (.CLK(clknet_leaf_272_clk_i),
    .D(_01903_),
    .Q(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _16765_ (.CLK(clknet_leaf_10_clk_i),
    .D(_01904_),
    .Q(\fifo0.fifo_store[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16766_ (.CLK(clknet_leaf_11_clk_i),
    .D(_01905_),
    .Q(\fifo0.fifo_store[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16767_ (.CLK(clknet_leaf_31_clk_i),
    .D(_01906_),
    .Q(\fifo0.fifo_store[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16768_ (.CLK(clknet_leaf_10_clk_i),
    .D(_01907_),
    .Q(\fifo0.fifo_store[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16769_ (.CLK(clknet_leaf_16_clk_i),
    .D(_01908_),
    .Q(\fifo0.fifo_store[79][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16770_ (.CLK(clknet_leaf_302_clk_i),
    .D(_01909_),
    .Q(\fifo0.fifo_store[79][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16771_ (.CLK(clknet_leaf_29_clk_i),
    .D(_01910_),
    .Q(\fifo0.fifo_store[79][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16772_ (.CLK(clknet_leaf_300_clk_i),
    .D(_01911_),
    .Q(\fifo0.fifo_store[79][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16773_ (.CLK(clknet_leaf_302_clk_i),
    .D(_01912_),
    .Q(\fifo0.fifo_store[79][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16774_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01913_),
    .Q(\fifo0.fifo_store[79][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16775_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01914_),
    .Q(\fifo0.fifo_store[79][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16776_ (.CLK(clknet_leaf_247_clk_i),
    .D(_01915_),
    .Q(\fifo0.fifo_store[79][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16777_ (.CLK(clknet_leaf_241_clk_i),
    .D(_01916_),
    .Q(\fifo0.fifo_store[79][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16778_ (.CLK(clknet_leaf_247_clk_i),
    .D(_01917_),
    .Q(\fifo0.fifo_store[79][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16779_ (.CLK(clknet_leaf_247_clk_i),
    .D(_01918_),
    .Q(\fifo0.fifo_store[79][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16780_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01919_),
    .Q(\fifo0.fifo_store[79][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16781_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01920_),
    .Q(\fifo0.fifo_store[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16782_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01921_),
    .Q(\fifo0.fifo_store[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16783_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01922_),
    .Q(\fifo0.fifo_store[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16784_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01923_),
    .Q(\fifo0.fifo_store[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16785_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01924_),
    .Q(\fifo0.fifo_store[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16786_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01925_),
    .Q(\fifo0.fifo_store[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16787_ (.CLK(clknet_leaf_331_clk_i),
    .D(_01926_),
    .Q(\fifo0.fifo_store[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16788_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01927_),
    .Q(\fifo0.fifo_store[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16789_ (.CLK(clknet_leaf_308_clk_i),
    .D(_01928_),
    .Q(\fifo0.fifo_store[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16790_ (.CLK(clknet_leaf_313_clk_i),
    .D(_01929_),
    .Q(\fifo0.fifo_store[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16791_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01930_),
    .Q(\fifo0.fifo_store[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16792_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01931_),
    .Q(\fifo0.fifo_store[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16793_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01932_),
    .Q(\fifo0.fifo_store[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16794_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01933_),
    .Q(\fifo0.fifo_store[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16795_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01934_),
    .Q(\fifo0.fifo_store[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16796_ (.CLK(clknet_leaf_274_clk_i),
    .D(_01935_),
    .Q(\fifo0.fifo_store[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16797_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01936_),
    .Q(\fifo0.fifo_store[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16798_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01937_),
    .Q(\fifo0.fifo_store[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16799_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01938_),
    .Q(\fifo0.fifo_store[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16800_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01939_),
    .Q(\fifo0.fifo_store[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16801_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01940_),
    .Q(\fifo0.fifo_store[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16802_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01941_),
    .Q(\fifo0.fifo_store[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16803_ (.CLK(clknet_leaf_310_clk_i),
    .D(_01942_),
    .Q(\fifo0.fifo_store[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16804_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01943_),
    .Q(\fifo0.fifo_store[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16805_ (.CLK(clknet_leaf_305_clk_i),
    .D(_01944_),
    .Q(\fifo0.fifo_store[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16806_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01945_),
    .Q(\fifo0.fifo_store[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16807_ (.CLK(clknet_leaf_267_clk_i),
    .D(_01946_),
    .Q(\fifo0.fifo_store[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16808_ (.CLK(clknet_leaf_254_clk_i),
    .D(_01947_),
    .Q(\fifo0.fifo_store[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16809_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01948_),
    .Q(\fifo0.fifo_store[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16810_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01949_),
    .Q(\fifo0.fifo_store[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16811_ (.CLK(clknet_leaf_256_clk_i),
    .D(_01950_),
    .Q(\fifo0.fifo_store[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16812_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01951_),
    .Q(\fifo0.fifo_store[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16813_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01952_),
    .Q(\fifo0.fifo_store[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16814_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01953_),
    .Q(\fifo0.fifo_store[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16815_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01954_),
    .Q(\fifo0.fifo_store[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16816_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01955_),
    .Q(\fifo0.fifo_store[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16817_ (.CLK(clknet_leaf_332_clk_i),
    .D(_01956_),
    .Q(\fifo0.fifo_store[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16818_ (.CLK(clknet_leaf_279_clk_i),
    .D(_01957_),
    .Q(\fifo0.fifo_store[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16819_ (.CLK(clknet_leaf_331_clk_i),
    .D(_01958_),
    .Q(\fifo0.fifo_store[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16820_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01959_),
    .Q(\fifo0.fifo_store[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16821_ (.CLK(clknet_leaf_307_clk_i),
    .D(_01960_),
    .Q(\fifo0.fifo_store[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16822_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01961_),
    .Q(\fifo0.fifo_store[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16823_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01962_),
    .Q(\fifo0.fifo_store[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16824_ (.CLK(clknet_leaf_270_clk_i),
    .D(_01963_),
    .Q(\fifo0.fifo_store[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16825_ (.CLK(clknet_leaf_263_clk_i),
    .D(_01964_),
    .Q(\fifo0.fifo_store[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16826_ (.CLK(clknet_leaf_261_clk_i),
    .D(_01965_),
    .Q(\fifo0.fifo_store[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16827_ (.CLK(clknet_leaf_262_clk_i),
    .D(_01966_),
    .Q(\fifo0.fifo_store[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16828_ (.CLK(clknet_leaf_274_clk_i),
    .D(_01967_),
    .Q(\fifo0.fifo_store[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16829_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01968_),
    .Q(\fifo0.fifo_store[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16830_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01969_),
    .Q(\fifo0.fifo_store[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16831_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01970_),
    .Q(\fifo0.fifo_store[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16832_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01971_),
    .Q(\fifo0.fifo_store[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16833_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01972_),
    .Q(\fifo0.fifo_store[127][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16834_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01973_),
    .Q(\fifo0.fifo_store[127][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16835_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01974_),
    .Q(\fifo0.fifo_store[127][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16836_ (.CLK(clknet_leaf_141_clk_i),
    .D(_01975_),
    .Q(\fifo0.fifo_store[127][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16837_ (.CLK(clknet_leaf_141_clk_i),
    .D(_01976_),
    .Q(\fifo0.fifo_store[127][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16838_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01977_),
    .Q(\fifo0.fifo_store[127][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16839_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01978_),
    .Q(\fifo0.fifo_store[127][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16840_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01979_),
    .Q(\fifo0.fifo_store[127][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16841_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01980_),
    .Q(\fifo0.fifo_store[127][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16842_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01981_),
    .Q(\fifo0.fifo_store[127][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16843_ (.CLK(clknet_leaf_175_clk_i),
    .D(_01982_),
    .Q(\fifo0.fifo_store[127][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16844_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01983_),
    .Q(\fifo0.fifo_store[127][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16845_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01984_),
    .Q(\dsmod0.mod2_ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16846_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01985_),
    .Q(\dsmod0.mod2_ctr[1] ));
 sky130_fd_sc_hd__dfxtp_4 _16847_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01986_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _16848_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01987_),
    .Q(\dsmod0.accu3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16849_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01988_),
    .Q(\dsmod0.accu3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16850_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01989_),
    .Q(\dsmod0.accu2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16851_ (.CLK(clknet_leaf_338_clk_i),
    .D(_01990_),
    .Q(\dsmod0.accu2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16852_ (.CLK(clknet_leaf_336_clk_i),
    .D(_01991_),
    .Q(\dsmod0.accu2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16853_ (.CLK(clknet_leaf_336_clk_i),
    .D(_01992_),
    .Q(\dsmod0.accu2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16854_ (.CLK(clknet_leaf_336_clk_i),
    .D(_01993_),
    .Q(\dsmod0.accu2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16855_ (.CLK(clknet_leaf_335_clk_i),
    .D(_01994_),
    .Q(\dsmod0.accu2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _16856_ (.CLK(clknet_leaf_335_clk_i),
    .D(_01995_),
    .Q(\dsmod0.accu2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16857_ (.CLK(clknet_leaf_329_clk_i),
    .D(_01996_),
    .Q(\dsmod0.accu2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _16858_ (.CLK(clknet_leaf_329_clk_i),
    .D(_01997_),
    .Q(\dsmod0.accu2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _16859_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01998_),
    .Q(\dsmod0.accu2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _16860_ (.CLK(clknet_leaf_327_clk_i),
    .D(_01999_),
    .Q(\dsmod0.accu2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _16861_ (.CLK(clknet_leaf_331_clk_i),
    .D(_02000_),
    .Q(\dsmod0.accu2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _16862_ (.CLK(clknet_leaf_331_clk_i),
    .D(_02001_),
    .Q(\dsmod0.accu2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _16863_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02002_),
    .Q(\dsmod0.accu2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _16864_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02003_),
    .Q(\dsmod0.accu2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _16865_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02004_),
    .Q(\dsmod0.accu2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _16866_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02005_),
    .Q(\dsmod0.accu1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16867_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02006_),
    .Q(\dsmod0.accu1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16868_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02007_),
    .Q(\dsmod0.accu1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16869_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02008_),
    .Q(\dsmod0.accu1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _16870_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02009_),
    .Q(\dsmod0.accu1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16871_ (.CLK(clknet_5_1_0_clk_i),
    .D(_02010_),
    .Q(\dsmod0.accu1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _16872_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02011_),
    .Q(\dsmod0.accu1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _16873_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02012_),
    .Q(\dsmod0.accu1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _16874_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02013_),
    .Q(\dsmod0.accu1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _16875_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02014_),
    .Q(\dsmod0.accu1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _16876_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02015_),
    .Q(\dsmod0.accu1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _16877_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02016_),
    .Q(\dsmod0.accu1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _16878_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02017_),
    .Q(\dsmod0.accu1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _16879_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02018_),
    .Q(\dsmod0.accu1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _16880_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02019_),
    .Q(\dsmod0.accu1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _16881_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02020_),
    .Q(\dsmod0.accu1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _16882_ (.CLK(clknet_leaf_2_clk_i),
    .D(_02021_),
    .Q(\fifo0.fifo_store[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16883_ (.CLK(clknet_leaf_4_clk_i),
    .D(_02022_),
    .Q(\fifo0.fifo_store[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16884_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02023_),
    .Q(\fifo0.fifo_store[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16885_ (.CLK(clknet_leaf_1_clk_i),
    .D(_02024_),
    .Q(\fifo0.fifo_store[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16886_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02025_),
    .Q(\fifo0.fifo_store[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16887_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02026_),
    .Q(\fifo0.fifo_store[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16888_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02027_),
    .Q(\fifo0.fifo_store[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16889_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02028_),
    .Q(\fifo0.fifo_store[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16890_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02029_),
    .Q(\fifo0.fifo_store[39][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16891_ (.CLK(clknet_leaf_22_clk_i),
    .D(_02030_),
    .Q(\fifo0.fifo_store[39][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16892_ (.CLK(clknet_leaf_290_clk_i),
    .D(_02031_),
    .Q(\fifo0.fifo_store[39][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16893_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02032_),
    .Q(\fifo0.fifo_store[39][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16894_ (.CLK(clknet_leaf_249_clk_i),
    .D(_02033_),
    .Q(\fifo0.fifo_store[39][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16895_ (.CLK(clknet_leaf_246_clk_i),
    .D(_02034_),
    .Q(\fifo0.fifo_store[39][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16896_ (.CLK(clknet_leaf_255_clk_i),
    .D(_02035_),
    .Q(\fifo0.fifo_store[39][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16897_ (.CLK(clknet_leaf_294_clk_i),
    .D(_02036_),
    .Q(\fifo0.fifo_store[39][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16898_ (.CLK(clknet_leaf_64_clk_i),
    .D(_02037_),
    .Q(\fifo0.fifo_store[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16899_ (.CLK(clknet_leaf_72_clk_i),
    .D(_02038_),
    .Q(\fifo0.fifo_store[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16900_ (.CLK(clknet_leaf_110_clk_i),
    .D(_02039_),
    .Q(\fifo0.fifo_store[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16901_ (.CLK(clknet_leaf_69_clk_i),
    .D(_02040_),
    .Q(\fifo0.fifo_store[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16902_ (.CLK(clknet_leaf_85_clk_i),
    .D(_02041_),
    .Q(\fifo0.fifo_store[119][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16903_ (.CLK(clknet_leaf_103_clk_i),
    .D(_02042_),
    .Q(\fifo0.fifo_store[119][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16904_ (.CLK(clknet_leaf_90_clk_i),
    .D(_02043_),
    .Q(\fifo0.fifo_store[119][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16905_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02044_),
    .Q(\fifo0.fifo_store[119][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16906_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02045_),
    .Q(\fifo0.fifo_store[119][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16907_ (.CLK(clknet_leaf_112_clk_i),
    .D(_02046_),
    .Q(\fifo0.fifo_store[119][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16908_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02047_),
    .Q(\fifo0.fifo_store[119][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16909_ (.CLK(clknet_leaf_178_clk_i),
    .D(_02048_),
    .Q(\fifo0.fifo_store[119][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16910_ (.CLK(clknet_leaf_178_clk_i),
    .D(_02049_),
    .Q(\fifo0.fifo_store[119][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16911_ (.CLK(clknet_leaf_160_clk_i),
    .D(_02050_),
    .Q(\fifo0.fifo_store[119][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16912_ (.CLK(clknet_leaf_178_clk_i),
    .D(_02051_),
    .Q(\fifo0.fifo_store[119][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16913_ (.CLK(clknet_leaf_158_clk_i),
    .D(_02052_),
    .Q(\fifo0.fifo_store[119][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16914_ (.CLK(clknet_leaf_62_clk_i),
    .D(_02053_),
    .Q(\fifo0.fifo_store[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16915_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02054_),
    .Q(\fifo0.fifo_store[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16916_ (.CLK(clknet_leaf_121_clk_i),
    .D(_02055_),
    .Q(\fifo0.fifo_store[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16917_ (.CLK(clknet_leaf_66_clk_i),
    .D(_02056_),
    .Q(\fifo0.fifo_store[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16918_ (.CLK(clknet_leaf_51_clk_i),
    .D(_02057_),
    .Q(\fifo0.fifo_store[69][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16919_ (.CLK(clknet_leaf_130_clk_i),
    .D(_02058_),
    .Q(\fifo0.fifo_store[69][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16920_ (.CLK(clknet_leaf_116_clk_i),
    .D(_02059_),
    .Q(\fifo0.fifo_store[69][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16921_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02060_),
    .Q(\fifo0.fifo_store[69][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16922_ (.CLK(clknet_leaf_127_clk_i),
    .D(_02061_),
    .Q(\fifo0.fifo_store[69][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16923_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02062_),
    .Q(\fifo0.fifo_store[69][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16924_ (.CLK(clknet_leaf_206_clk_i),
    .D(_02063_),
    .Q(\fifo0.fifo_store[69][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16925_ (.CLK(clknet_leaf_198_clk_i),
    .D(_02064_),
    .Q(\fifo0.fifo_store[69][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16926_ (.CLK(clknet_leaf_201_clk_i),
    .D(_02065_),
    .Q(\fifo0.fifo_store[69][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16927_ (.CLK(clknet_leaf_201_clk_i),
    .D(_02066_),
    .Q(\fifo0.fifo_store[69][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16928_ (.CLK(clknet_leaf_199_clk_i),
    .D(_02067_),
    .Q(\fifo0.fifo_store[69][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16929_ (.CLK(clknet_leaf_207_clk_i),
    .D(_02068_),
    .Q(\fifo0.fifo_store[69][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16930_ (.CLK(clknet_leaf_328_clk_i),
    .D(_02069_),
    .Q(\dsmod0.mod2_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16931_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02070_),
    .Q(\dsmod0.mod2_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _16932_ (.CLK(clknet_leaf_56_clk_i),
    .D(_02071_),
    .Q(\fifo0.fifo_store[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16933_ (.CLK(clknet_leaf_12_clk_i),
    .D(_02072_),
    .Q(\fifo0.fifo_store[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16934_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02073_),
    .Q(\fifo0.fifo_store[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16935_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02074_),
    .Q(\fifo0.fifo_store[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16936_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02075_),
    .Q(\fifo0.fifo_store[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16937_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02076_),
    .Q(\fifo0.fifo_store[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16938_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02077_),
    .Q(\fifo0.fifo_store[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16939_ (.CLK(clknet_leaf_215_clk_i),
    .D(_02078_),
    .Q(\fifo0.fifo_store[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16940_ (.CLK(clknet_leaf_33_clk_i),
    .D(_02079_),
    .Q(\fifo0.fifo_store[47][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16941_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02080_),
    .Q(\fifo0.fifo_store[47][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16942_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02081_),
    .Q(\fifo0.fifo_store[47][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16943_ (.CLK(clknet_leaf_249_clk_i),
    .D(_02082_),
    .Q(\fifo0.fifo_store[47][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16944_ (.CLK(clknet_leaf_240_clk_i),
    .D(_02083_),
    .Q(\fifo0.fifo_store[47][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16945_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02084_),
    .Q(\fifo0.fifo_store[47][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16946_ (.CLK(clknet_leaf_239_clk_i),
    .D(_02085_),
    .Q(\fifo0.fifo_store[47][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16947_ (.CLK(clknet_leaf_293_clk_i),
    .D(_02086_),
    .Q(\fifo0.fifo_store[47][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16948_ (.CLK(clknet_leaf_2_clk_i),
    .D(_02087_),
    .Q(\fifo0.fifo_store[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16949_ (.CLK(clknet_leaf_3_clk_i),
    .D(_02088_),
    .Q(\fifo0.fifo_store[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16950_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02089_),
    .Q(\fifo0.fifo_store[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16951_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02090_),
    .Q(\fifo0.fifo_store[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16952_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02091_),
    .Q(\fifo0.fifo_store[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16953_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02092_),
    .Q(\fifo0.fifo_store[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16954_ (.CLK(clknet_leaf_317_clk_i),
    .D(_02093_),
    .Q(\fifo0.fifo_store[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16955_ (.CLK(clknet_leaf_284_clk_i),
    .D(_02094_),
    .Q(\fifo0.fifo_store[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16956_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02095_),
    .Q(\fifo0.fifo_store[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16957_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02096_),
    .Q(\fifo0.fifo_store[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16958_ (.CLK(clknet_leaf_268_clk_i),
    .D(_02097_),
    .Q(\fifo0.fifo_store[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16959_ (.CLK(clknet_leaf_267_clk_i),
    .D(_02098_),
    .Q(\fifo0.fifo_store[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16960_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02099_),
    .Q(\fifo0.fifo_store[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16961_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02100_),
    .Q(\fifo0.fifo_store[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16962_ (.CLK(clknet_leaf_263_clk_i),
    .D(_02101_),
    .Q(\fifo0.fifo_store[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16963_ (.CLK(clknet_leaf_286_clk_i),
    .D(_02102_),
    .Q(\fifo0.fifo_store[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16964_ (.CLK(clknet_leaf_63_clk_i),
    .D(_02103_),
    .Q(\fifo0.fifo_store[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16965_ (.CLK(clknet_leaf_73_clk_i),
    .D(_02104_),
    .Q(\fifo0.fifo_store[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16966_ (.CLK(clknet_leaf_117_clk_i),
    .D(_02105_),
    .Q(\fifo0.fifo_store[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16967_ (.CLK(clknet_leaf_67_clk_i),
    .D(_02106_),
    .Q(\fifo0.fifo_store[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16968_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02107_),
    .Q(\fifo0.fifo_store[109][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16969_ (.CLK(clknet_leaf_108_clk_i),
    .D(_02108_),
    .Q(\fifo0.fifo_store[109][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16970_ (.CLK(clknet_leaf_115_clk_i),
    .D(_02109_),
    .Q(\fifo0.fifo_store[109][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16971_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02110_),
    .Q(\fifo0.fifo_store[109][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16972_ (.CLK(clknet_leaf_118_clk_i),
    .D(_02111_),
    .Q(\fifo0.fifo_store[109][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16973_ (.CLK(clknet_leaf_113_clk_i),
    .D(_02112_),
    .Q(\fifo0.fifo_store[109][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16974_ (.CLK(clknet_leaf_160_clk_i),
    .D(_02113_),
    .Q(\fifo0.fifo_store[109][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16975_ (.CLK(clknet_leaf_177_clk_i),
    .D(_02114_),
    .Q(\fifo0.fifo_store[109][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16976_ (.CLK(clknet_leaf_173_clk_i),
    .D(_02115_),
    .Q(\fifo0.fifo_store[109][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16977_ (.CLK(clknet_leaf_176_clk_i),
    .D(_02116_),
    .Q(\fifo0.fifo_store[109][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16978_ (.CLK(clknet_leaf_183_clk_i),
    .D(_02117_),
    .Q(\fifo0.fifo_store[109][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16979_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02118_),
    .Q(\fifo0.fifo_store[109][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16980_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02119_),
    .Q(\sinegen0.read_ptr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _16981_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02120_),
    .Q(\sinegen0.read_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16982_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02121_),
    .Q(\sinegen0.read_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16983_ (.CLK(clknet_leaf_5_clk_i),
    .D(_02122_),
    .Q(\sinegen0.read_ptr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _16984_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02123_),
    .Q(\sinegen0.read_ptr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _16985_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02124_),
    .Q(\sinegen0.read_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _16986_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02125_),
    .Q(\sinegen0.read_ptr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16987_ (.CLK(clknet_leaf_57_clk_i),
    .D(_02126_),
    .Q(\fifo0.fifo_store[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16988_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02127_),
    .Q(\fifo0.fifo_store[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16989_ (.CLK(clknet_leaf_115_clk_i),
    .D(_02128_),
    .Q(\fifo0.fifo_store[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16990_ (.CLK(clknet_leaf_49_clk_i),
    .D(_02129_),
    .Q(\fifo0.fifo_store[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16991_ (.CLK(clknet_leaf_52_clk_i),
    .D(_02130_),
    .Q(\fifo0.fifo_store[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16992_ (.CLK(clknet_leaf_119_clk_i),
    .D(_02131_),
    .Q(\fifo0.fifo_store[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16993_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02132_),
    .Q(\fifo0.fifo_store[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16994_ (.CLK(clknet_leaf_128_clk_i),
    .D(_02133_),
    .Q(\fifo0.fifo_store[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16995_ (.CLK(clknet_leaf_122_clk_i),
    .D(_02134_),
    .Q(\fifo0.fifo_store[50][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16996_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02135_),
    .Q(\fifo0.fifo_store[50][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16997_ (.CLK(clknet_leaf_223_clk_i),
    .D(_02136_),
    .Q(\fifo0.fifo_store[50][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16998_ (.CLK(clknet_leaf_196_clk_i),
    .D(_02137_),
    .Q(\fifo0.fifo_store[50][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16999_ (.CLK(clknet_leaf_235_clk_i),
    .D(_02138_),
    .Q(\fifo0.fifo_store[50][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17000_ (.CLK(clknet_leaf_195_clk_i),
    .D(_02139_),
    .Q(\fifo0.fifo_store[50][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17001_ (.CLK(clknet_leaf_234_clk_i),
    .D(_02140_),
    .Q(\fifo0.fifo_store[50][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17002_ (.CLK(clknet_leaf_221_clk_i),
    .D(_02141_),
    .Q(\fifo0.fifo_store[50][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17003_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02142_),
    .Q(\fifo0.fifo_store[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17004_ (.CLK(clknet_leaf_78_clk_i),
    .D(_02143_),
    .Q(\fifo0.fifo_store[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17005_ (.CLK(clknet_leaf_91_clk_i),
    .D(_02144_),
    .Q(\fifo0.fifo_store[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17006_ (.CLK(clknet_leaf_68_clk_i),
    .D(_02145_),
    .Q(\fifo0.fifo_store[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17007_ (.CLK(clknet_leaf_85_clk_i),
    .D(_02146_),
    .Q(\fifo0.fifo_store[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17008_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02147_),
    .Q(\fifo0.fifo_store[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17009_ (.CLK(clknet_leaf_97_clk_i),
    .D(_02148_),
    .Q(\fifo0.fifo_store[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17010_ (.CLK(clknet_leaf_215_clk_i),
    .D(_02149_),
    .Q(\fifo0.fifo_store[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17011_ (.CLK(clknet_leaf_33_clk_i),
    .D(_02150_),
    .Q(\fifo0.fifo_store[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17012_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02151_),
    .Q(\fifo0.fifo_store[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17013_ (.CLK(clknet_leaf_198_clk_i),
    .D(_02152_),
    .Q(\fifo0.fifo_store[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17014_ (.CLK(clknet_leaf_200_clk_i),
    .D(_02153_),
    .Q(\fifo0.fifo_store[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17015_ (.CLK(clknet_leaf_193_clk_i),
    .D(_02154_),
    .Q(\fifo0.fifo_store[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17016_ (.CLK(clknet_leaf_187_clk_i),
    .D(_02155_),
    .Q(\fifo0.fifo_store[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17017_ (.CLK(clknet_leaf_188_clk_i),
    .D(_02156_),
    .Q(\fifo0.fifo_store[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17018_ (.CLK(clknet_leaf_207_clk_i),
    .D(_02157_),
    .Q(\fifo0.fifo_store[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17019_ (.CLK(clknet_leaf_279_clk_i),
    .D(_02158_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_1 _17020_ (.CLK(clknet_leaf_279_clk_i),
    .D(_02159_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_4 _17021_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02160_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_2 _17022_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02161_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_4 _17023_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02162_),
    .Q(_00004_));
 sky130_fd_sc_hd__dfxtp_4 _17024_ (.CLK(clknet_leaf_277_clk_i),
    .D(_02163_),
    .Q(_00005_));
 sky130_fd_sc_hd__dfxtp_4 _17025_ (.CLK(clknet_leaf_277_clk_i),
    .D(_02164_),
    .Q(_00006_));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(fifo_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(fifo_i[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(fifo_i[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(fifo_i[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(fifo_i[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(fifo_i[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(fifo_i[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(fifo_i[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(fifo_i[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(fifo_i[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(fifo_i[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(fifo_i[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(fifo_i[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(fifo_i[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(fifo_i[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(fifo_i[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(fifo_rdy_i),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(mode_i),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(osr_i[0]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(osr_i[1]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(rst_n_i),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(tst_fifo_loop_i),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(tst_sinegen_en_i),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(tst_sinegen_step_i[0]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(tst_sinegen_step_i[1]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(tst_sinegen_step_i[2]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(tst_sinegen_step_i[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(tst_sinegen_step_i[4]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(tst_sinegen_step_i[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(volume_i[0]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(volume_i[1]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(volume_i[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(volume_i[3]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(ds_n_o));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(ds_o));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(fifo_ack_o));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(fifo_empty_o));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(fifo_full_o));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_5_2_0_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_5_3_0_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i (.A(clknet_5_8_0_clk_i),
    .X(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i (.A(clknet_5_9_0_clk_i),
    .X(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i (.A(clknet_5_10_0_clk_i),
    .X(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i (.A(clknet_5_11_0_clk_i),
    .X(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_108_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk_i (.A(clknet_5_15_0_clk_i),
    .X(clknet_leaf_109_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_110_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_111_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk_i (.A(clknet_5_14_0_clk_i),
    .X(clknet_leaf_112_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_113_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_114_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk_i (.A(clknet_5_12_0_clk_i),
    .X(clknet_leaf_115_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_116_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_117_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_118_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_119_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_120_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_121_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_122_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_123_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk_i (.A(clknet_5_13_0_clk_i),
    .X(clknet_leaf_124_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_125_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_126_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_127_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_128_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_129_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_130_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_131_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_132_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_133_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_134_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_135_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_136_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_137_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_138_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_139_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_140_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_141_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_142_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_143_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_144_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_145_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_146_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_147_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_148_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_149_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_150_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk_i (.A(clknet_5_26_0_clk_i),
    .X(clknet_leaf_151_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_152_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_153_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_154_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_155_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_156_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_157_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_158_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk_i (.A(clknet_5_27_0_clk_i),
    .X(clknet_leaf_159_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_160_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_161_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_162_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_163_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_164_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_165_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_166_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_167_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_168_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_169_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_170_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_171_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_172_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_173_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_174_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk_i (.A(clknet_5_31_0_clk_i),
    .X(clknet_leaf_175_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_176_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_177_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_178_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_179_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_180_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_181_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_182_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_183_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_184_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_185_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_186_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_187_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_188_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_189_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_190_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_191_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk_i (.A(clknet_5_29_0_clk_i),
    .X(clknet_leaf_192_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_193_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_194_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_195_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_196_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_197_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_198_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_199_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_200_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_201_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_202_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_203_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk_i (.A(clknet_5_30_0_clk_i),
    .X(clknet_leaf_204_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_205_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_206_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_207_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_208_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk_i (.A(clknet_5_28_0_clk_i),
    .X(clknet_leaf_209_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_210_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_211_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk_i (.A(clknet_5_25_0_clk_i),
    .X(clknet_leaf_212_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_213_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_214_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_215_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk_i (.A(clknet_5_24_0_clk_i),
    .X(clknet_leaf_216_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_217_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_218_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_219_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_220_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_221_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_222_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_223_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_224_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_225_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_226_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_227_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_228_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_229_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_230_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_231_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_232_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_233_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk_i (.A(clknet_5_22_0_clk_i),
    .X(clknet_leaf_234_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_235_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_236_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_237_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_238_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_239_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_240_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_241_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_242_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_243_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_244_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_245_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_246_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_247_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk_i (.A(clknet_5_23_0_clk_i),
    .X(clknet_leaf_248_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_249_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_250_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_251_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_252_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_253_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_254_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_255_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_256_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_257_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk_i (.A(clknet_5_21_0_clk_i),
    .X(clknet_leaf_258_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_259_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_260_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_261_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_262_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_263_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_264_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk_i (.A(clknet_5_20_0_clk_i),
    .X(clknet_leaf_265_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_266_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_267_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_268_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_269_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_270_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_271_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_272_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_273_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_274_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_275_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_277_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_278_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_279_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_280_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_281_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_282_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_283_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_284_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk_i (.A(clknet_5_16_0_clk_i),
    .X(clknet_leaf_285_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_286_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_287_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_288_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk_i (.A(clknet_5_17_0_clk_i),
    .X(clknet_leaf_289_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_290_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_291_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_292_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_293_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk_i (.A(clknet_5_19_0_clk_i),
    .X(clknet_leaf_294_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_295_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_296_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_297_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_298_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_299_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_300_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_clk_i (.A(clknet_5_18_0_clk_i),
    .X(clknet_leaf_301_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_302_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_303_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_304_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_305_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_306_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_306_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_307_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_308_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_309_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_clk_i (.A(clknet_5_7_0_clk_i),
    .X(clknet_leaf_310_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_311_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_312_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_clk_i (.A(clknet_5_6_0_clk_i),
    .X(clknet_leaf_313_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_314_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_315_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_316_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_317_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_318_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_319_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_320_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_321_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_322_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_323_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_324_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_324_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_clk_i (.A(clknet_5_5_0_clk_i),
    .X(clknet_leaf_325_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_326_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_326_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_327_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_328_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_329_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_330_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_331_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_clk_i (.A(clknet_5_4_0_clk_i),
    .X(clknet_leaf_332_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_333_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_333_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_335_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_335_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_336_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_336_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_337_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_337_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_338_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_338_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_339_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_339_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_340_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_340_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_341_clk_i (.A(clknet_5_0_0_clk_i),
    .X(clknet_leaf_341_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_342_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_342_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_343_clk_i (.A(clknet_5_1_0_clk_i),
    .X(clknet_leaf_343_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_clk_i (.A(clknet_1_0_0_clk_i),
    .X(clknet_1_0_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_clk_i (.A(clknet_1_1_0_clk_i),
    .X(clknet_1_1_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk_i (.A(clknet_1_0_1_clk_i),
    .X(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_1_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_2_0_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk_i (.A(clknet_1_0_1_clk_i),
    .X(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_1_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_2_1_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk_i (.A(clknet_1_1_1_clk_i),
    .X(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_1_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_2_2_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk_i (.A(clknet_1_1_1_clk_i),
    .X(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_1_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_2_3_1_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk_i (.A(clknet_2_0_1_clk_i),
    .X(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk_i (.A(clknet_2_0_1_clk_i),
    .X(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk_i (.A(clknet_2_1_1_clk_i),
    .X(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk_i (.A(clknet_2_1_1_clk_i),
    .X(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk_i (.A(clknet_2_2_1_clk_i),
    .X(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk_i (.A(clknet_2_2_1_clk_i),
    .X(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk_i (.A(clknet_2_3_1_clk_i),
    .X(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk_i (.A(clknet_2_3_1_clk_i),
    .X(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk_i (.A(clknet_3_0_0_clk_i),
    .X(clknet_4_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk_i (.A(clknet_3_0_0_clk_i),
    .X(clknet_4_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk_i (.A(clknet_3_1_0_clk_i),
    .X(clknet_4_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk_i (.A(clknet_3_1_0_clk_i),
    .X(clknet_4_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk_i (.A(clknet_3_2_0_clk_i),
    .X(clknet_4_4_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk_i (.A(clknet_3_2_0_clk_i),
    .X(clknet_4_5_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk_i (.A(clknet_3_3_0_clk_i),
    .X(clknet_4_6_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk_i (.A(clknet_3_3_0_clk_i),
    .X(clknet_4_7_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk_i (.A(clknet_3_4_0_clk_i),
    .X(clknet_4_8_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk_i (.A(clknet_3_4_0_clk_i),
    .X(clknet_4_9_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk_i (.A(clknet_3_5_0_clk_i),
    .X(clknet_4_10_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk_i (.A(clknet_3_5_0_clk_i),
    .X(clknet_4_11_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk_i (.A(clknet_3_6_0_clk_i),
    .X(clknet_4_12_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk_i (.A(clknet_3_6_0_clk_i),
    .X(clknet_4_13_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk_i (.A(clknet_3_7_0_clk_i),
    .X(clknet_4_14_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk_i (.A(clknet_3_7_0_clk_i),
    .X(clknet_4_15_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_0_0_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_1_0_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_2_0_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_3_0_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_4_0_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_5_0_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_6_0_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_7_0_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_8_0_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_9_0_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_10_0_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_11_0_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_12_0_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_13_0_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_14_0_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_15_0_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_16_0_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_17_0_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_18_0_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_19_0_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_20_0_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_21_0_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_22_0_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_23_0_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_24_0_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_25_0_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_26_0_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_27_0_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_28_0_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_29_0_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_30_0_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_31_0_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__C1 (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__B1 (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__B1 (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__A (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__B1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__B1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__C1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__B1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__B (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__A (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__C (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__B (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A2 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__B1 (.DIODE(_02192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13886__A (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13369__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__A2 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14111__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__A (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A1 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A2 (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__S0 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__S0 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13470__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__A1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__A_N (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13331__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__B2 (.DIODE(_02270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A2 (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A2 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__C1 (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A3 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13517__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13327__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__A2 (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__C1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__C1 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A2 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__B1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__B1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A3 (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A2 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__C1 (.DIODE(_02537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__A2 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__B1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A3 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__B2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__B1 (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__C1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__B (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__A2 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__B1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__B (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A2 (.DIODE(_02606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A2 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__B1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A2 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A2 (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__B1 (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__A2 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__A1 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__A2 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13567__B (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__B2 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A3 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A2 (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__B1 (.DIODE(_02692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13614__A1 (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__B1 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__B1 (.DIODE(_02701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A2 (.DIODE(_02708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__B1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__B (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__A0 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__A2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__B1 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A3 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A2 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__C1 (.DIODE(_02791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13729__B1 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__B (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__A2 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__B (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__B (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__A2 (.DIODE(_02836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__B (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__B (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__B2 (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__A2 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__A2 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__A2 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14143__A1 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__B_N (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14114__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14078__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13808__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13783__S0 (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14114__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14078__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13808__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13793__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13783__S1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14145__C1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__A (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14118__A (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14113__B1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14093__A1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__A (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__B1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__A1 (.DIODE(_02866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14146__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14131__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__S0 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A2 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14112__S (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14096__S (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14063__S0 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14052__S0 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__S0 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14000__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13887__A1 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__S (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__S (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13793__A2 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__B1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14129__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14106__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14080__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__S0 (.DIODE(_02878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14129__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14071__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__S1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__A2 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14147__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14136__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14126__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14057__B1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__S1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__S1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__S1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__C1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14011__B1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__S1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__C1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__S1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13817__A (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A2 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__B (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__B2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13885__A1 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13877__A1 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13841__A2 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13870__A2 (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__B1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__C1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__B (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A2 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__A2 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13908__A2 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14049__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14047__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14038__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14008__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__S1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__A (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A2 (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__A0 (.DIODE(_02999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__B2 (.DIODE(_03005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__B1 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A1_N (.DIODE(_03008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13935__B (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A1 (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__C1 (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__B1 (.DIODE(_03035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13955__A2 (.DIODE(_03036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13963__A2 (.DIODE(_03044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A2_N (.DIODE(_03048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__A1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14132__A1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14124__A (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__A1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__A1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__C1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14050__A (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__C1 (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__A (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__A1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__A1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__A (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__A (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__B1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__A1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__B1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A1 (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14057__A1 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__S0 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__S0 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__S (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14028__A (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14011__A1 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__S0 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__S (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__S0 (.DIODE(_03063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14061__A (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__A (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14044__A1 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__A1 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__B2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A1 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14009__A (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__B2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__A (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14049__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14047__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14038__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14008__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__S0 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14044__B1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__B1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__C1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__C1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__C1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__C1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14006__A1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__C1 (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__S (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__S (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14002__S0 (.DIODE(_03082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14111__C1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__C1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14002__S1 (.DIODE(_03083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__B (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__A3 (.DIODE(_03119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14040__A0 (.DIODE(_03120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__A2 (.DIODE(_03122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__A2 (.DIODE(_03130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__B (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__B2 (.DIODE(_03149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__A2 (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__B (.DIODE(_03153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__B1 (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__B (.DIODE(_03162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14109__A2 (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A2 (.DIODE(_03185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__A2 (.DIODE(_03198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14118__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14122__A0 (.DIODE(_03202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__B1 (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14130__B (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14136__A2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14139__B (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14147__A2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__B2 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14160__A2 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14151__B (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14222__A2 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14213__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__B (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__B (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14227__B (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14226__B (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__B1 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__B1 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__A1 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14255__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__B2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__A1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__A (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__B2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__B2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14371__A (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__A1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__B2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14245__A2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__A1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14502__B1 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__B1 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__A1 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14386__A (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__A (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__A1 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__B (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__B (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__A (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__A (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14274__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14270__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14264__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14262__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14260__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__A2 (.DIODE(_03328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14647__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__B (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14265__B (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14252__B (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14274__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14270__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14264__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14262__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14260__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__C1 (.DIODE(_03332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14645__A2_N (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14344__B2 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14263__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14261__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14259__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__B (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14375__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14345__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14329__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14533__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14466__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14403__C1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14375__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14345__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14329__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14299__A2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__B1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__A (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__C1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A2_N (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14487__B2 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__C1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__B1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__A2 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__C1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__B1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__B (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14296__B1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14779__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14647__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14533__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14466__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14299__C1 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14560__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__S (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__A (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14554__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14540__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14538__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__S (.DIODE(_03582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14600__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14569__A (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14582__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14578__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14576__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__S (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14630__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14628__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__S (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14603__A (.DIODE(_03617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14620__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14618__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14612__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14678__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14670__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__A (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14660__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14654__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__S (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14708__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14706__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__S (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14683__A (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14702__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14700__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14696__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14694__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14690__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14744__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14742__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14740__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14738__S (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__A (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14736__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14734__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14730__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14724__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14722__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14720__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14718__S (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14779__A2 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14778__A (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A2 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14771__A (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__A2 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14764__A (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__A2 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__B1 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14753__A3 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__A2 (.DIODE(_03700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__A2 (.DIODE(_03721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14777__B (.DIODE(_03721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14821__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14819__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__S (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14794__A (.DIODE(_03735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14811__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14801__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14795__S (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14859__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14853__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14849__S (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__A (.DIODE(_03753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14845__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14841__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14839__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14835__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14829__S (.DIODE(_03754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A2 (.DIODE(_03779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(_03779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__B1 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A1 (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(_03814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A2 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__B (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B2 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__B2 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__B2 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B2 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__B (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A0 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14829__A1 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09069__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A0 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A2 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A2 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A1 (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__C (.DIODE(_03824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__A2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A2 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B1 (.DIODE(_03827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A0 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__B1 (.DIODE(_03829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__B2 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A0 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B1 (.DIODE(_03832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A0 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B1 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A0 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A (.DIODE(_03837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A (.DIODE(_03837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A (.DIODE(_03838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A0 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B1 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A0 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B1 (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__A0 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B1 (.DIODE(_03844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A0 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B1 (.DIODE(_03846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A0 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B1 (.DIODE(_03848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A (.DIODE(_03849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A (.DIODE(_03849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(_03850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A0 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__B1 (.DIODE(_03851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__A0 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B1 (.DIODE(_03854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A0 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__B1 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A0 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__B1 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A0 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B1 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__A (.DIODE(_03861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(_03861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A (.DIODE(_03861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A (.DIODE(_03861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A0 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A3 (.DIODE(_03862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A (.DIODE(_03866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__B (.DIODE(_03866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A (.DIODE(_03866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__B (.DIODE(_03866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__S (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__A1 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A (.DIODE(_03875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A1 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14839__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14694__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14660__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14618__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A1 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A (.DIODE(_03896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(_03897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14849__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14738__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14670__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A1 (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__A (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A1 (.DIODE(_03900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14740__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14706__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A1 (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A (.DIODE(_03902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A1 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14853__A1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14819__A1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__A1 (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A (.DIODE(_03908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A1 (.DIODE(_03909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__A1 (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08643__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A (.DIODE(_03911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A1 (.DIODE(_03912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14859__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A1 (.DIODE(_03915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14648__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14568__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A (.DIODE(_03919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__B (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__S (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__A (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__S (.DIODE(_03922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__B (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__B (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__S (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__S (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14682__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14602__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__B (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__B (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__B (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__S (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(_03966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__S (.DIODE(_03967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__A (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__B (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__B (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__B (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__B (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__B (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__A (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A (.DIODE(_03986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14793__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A (.DIODE(_03989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__B (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__B (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__S (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A (.DIODE(_03991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__S (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__A (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__B (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__S (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__S (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A (.DIODE(_04031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__B (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__B (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__S (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__B (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__B (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__S (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__S (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__S (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__S (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__S (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__S (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__S (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__S (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__S (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14602__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__B (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__S (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__S (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A1 (.DIODE(_04153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__A1 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__B (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__B (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__B (.DIODE(_04172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__S (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__A (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__S (.DIODE(_04174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08575__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A1 (.DIODE(_04182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A1 (.DIODE(_04190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A1 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(_04199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__S (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__S (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__A (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__S (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__S (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__S (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A (.DIODE(_04259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__B (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__B (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__S (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__S (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__B (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__S (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A (.DIODE(_04298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__S (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14568__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__S (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(_04319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__S (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A (.DIODE(_04337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__S (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__S (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__S (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__B (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__S (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A (.DIODE(_04377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__S (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__S (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__S (.DIODE(_04396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__S (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__A (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__S (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__S (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__S (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A1 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__A1 (.DIODE(_04441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__S (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08575__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__S (.DIODE(_04454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A1 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__S (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__A (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__S (.DIODE(_04474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A1 (.DIODE(_04476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__A1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A1 (.DIODE(_04482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A1 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A1 (.DIODE(_04488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A1 (.DIODE(_04494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A1 (.DIODE(_04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__S (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__S (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__S (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__S (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__A (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__S (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__S (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__S (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__S (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__S (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__S (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__S (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__S (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__S (.DIODE(_04632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__S (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__S (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A1 (.DIODE(_04656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09015__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A1 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A1 (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__S (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__S (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__S (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__A (.DIODE(_04691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09015__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__S (.DIODE(_04692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__A1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__S (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A (.DIODE(_04730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A1 (.DIODE(_04733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A1 (.DIODE(_04735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A1 (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A1 (.DIODE(_04739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A1 (.DIODE(_04742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A1 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__A1 (.DIODE(_04751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__S (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__S (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A (.DIODE(_04794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__S (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__S (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__S (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__S (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__S (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09320__A (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__S (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A0 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__S (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A (.DIODE(_04887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__S (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A0 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A0 (.DIODE(_04892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A0 (.DIODE(_04894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A0 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A0 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A0 (.DIODE(_04900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A0 (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A0 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A0 (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A0 (.DIODE(_04910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A0 (.DIODE(_04912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A0 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A0 (.DIODE(_04916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A0 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__A (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A1 (.DIODE(_04927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A1 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__S (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__S (.DIODE(_04943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__S (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__S (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__S (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(_04981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__A1 (.DIODE(_04997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A1 (.DIODE(_04999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B (.DIODE(_05001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__S (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__S (.DIODE(_05003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__A1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__S (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__S (.DIODE(_05048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__A (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__A (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__S (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__A (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__S (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__S (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__A (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A1 (.DIODE(_05153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__S (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__S (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__S (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__A (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__S (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__S (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__S (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__A1 (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__S (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__S (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__S (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__A (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__A1 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__A1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__A1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A1 (.DIODE(_05256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__A1 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__S (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__S (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__S (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__S (.DIODE(_05282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__S (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__S (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__S (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__S (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__S (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__S (.DIODE(_05337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__S (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__A (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__S (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__S (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A (.DIODE(_05372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__S (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__S (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A1 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A1 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A1 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A1 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__S (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(_05412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__S (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__S (.DIODE(_05431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__S (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__A (.DIODE(_05449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__S (.DIODE(_05450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__S (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__S (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A1 (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A1 (.DIODE(_05486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A1 (.DIODE(_05488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__S (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__S (.DIODE(_05490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__A1 (.DIODE(_05503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A1 (.DIODE(_05505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__S (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__S (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__S (.DIODE(_05534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__S (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__S (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__S (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__S (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__S (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A (.DIODE(_05590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__S (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__S (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A (.DIODE(_05608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__S (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__S (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__S (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__S (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A (.DIODE(_05645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__S (.DIODE(_05646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A1 (.DIODE(_05652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__A1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__A1 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__S (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__S (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__S (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__S (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__S (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__A1 (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__S (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__A (.DIODE(_05722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__S (.DIODE(_05723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A1 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A1 (.DIODE(_05741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__S (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A (.DIODE(_05743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__S (.DIODE(_05744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__S (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A (.DIODE(_05762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__S (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A1 (.DIODE(_05768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A1 (.DIODE(_05770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__S (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__S (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__S (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__S (.DIODE(_05809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__S (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__A (.DIODE(_05826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__S (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__S (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__S (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__S (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A (.DIODE(_05862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__S (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(_05872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A1 (.DIODE(_05876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11341__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A1 (.DIODE(_05878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__S (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__C1 (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14298__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14277__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14238__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__B1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__C1 (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A (.DIODE(_05903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14753__C1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__A (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14520__B1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14453__B1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14246__A (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__B1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B1 (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A (.DIODE(_05924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14423__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14358__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__C1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__B1 (.DIODE(_05927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__C (.DIODE(_05943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A2 (.DIODE(_05943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B (.DIODE(_05943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__S (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11341__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__S (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__S (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__S (.DIODE(_05997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11418__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__S (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A (.DIODE(_06014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__S (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A1 (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A1 (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__S (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A (.DIODE(_06034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__S (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__A1 (.DIODE(_06037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A1 (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__S (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A1 (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A1 (.DIODE(_06061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A1 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A1 (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__S (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(_06080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__S (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__S (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__A (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__S (.DIODE(_06099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__S (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__S (.DIODE(_06117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A1 (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A1 (.DIODE(_06126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__A1 (.DIODE(_06130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A1 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__S (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__A (.DIODE(_06138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__S (.DIODE(_06139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__S (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__S (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__S (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__S (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__S (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__A (.DIODE(_06232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__S (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__S (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11872__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__S (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__S (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14742__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14708__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14628__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14560__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11872__A1 (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14795__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14718__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A1 (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__S (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__S (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14720__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14538__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A1 (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14821__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14744__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14630__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14678__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A1 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14600__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A1 (.DIODE(_06304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__S (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11929__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__S (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14722__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14654__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14540__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__A1 (.DIODE(_06310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14835__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14801__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14724__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14690__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14576__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11929__A1 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14612__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14578__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A1 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14841__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14730__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14696__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14582__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__A1 (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14845__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14811__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14734__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14700__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14620__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14736__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14702__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14554__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11960__A (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__S (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__B2 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__B1 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14462__B1 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14441__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14343__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14293__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__B1 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__B1 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14504__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14432__B1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14403__B2 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14344__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14328__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A2 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14164__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__B1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13975__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__C1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__C (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A1 (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__C (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__A1 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14225__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__C1 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__B1 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__B1 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__B1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__B1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__B1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__B1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__C1 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13667__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13575__B1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__C1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__S (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__B1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14779__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14773__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__C1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__B1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__C1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__B (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__B (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A2 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A1 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__B (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A2 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A2 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A2 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A2 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__B1 (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__B1 (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A1 (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12415__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A (.DIODE(_06362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13575__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__C1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__B1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A1 (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__A (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__C1 (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__C1 (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__S0 (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A1 (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__A1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__C1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13286__A1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__B1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__B1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__C1 (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13967__A1 (.DIODE(_06374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13282__C1 (.DIODE(_06374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__B (.DIODE(_06374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__B (.DIODE(_06374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__B1_N (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__B1_N (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__A_N (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__B1 (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__B1 (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13674__A1 (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__A (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__C1 (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__A1 (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__A1 (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__C1 (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__A (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A (.DIODE(_06377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__A (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__B1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__A1 (.DIODE(_06378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14759__A1 (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__A1 (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__A (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__C1 (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__C (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__B (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A2 (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__B (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__C (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__A (.DIODE(_06380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A2 (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A2 (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__B (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A2 (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__A3 (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__B2 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A2 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A1 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__C1 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A1 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A2 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__B1 (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__A (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__A1 (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__B (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__B (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__A1 (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A1 (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__B (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12415__C_N (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__A (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__B1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__B1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__A1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__B1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13667__A1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13574__B1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__A (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__A1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__B1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__B1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A1 (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__A (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__B1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__A1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__B1 (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A (.DIODE(_06397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__A1 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14761__A (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14760__A (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A2 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A1 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A1 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__A1 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__B (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__A1 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__A (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14753__A1 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__B1 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__B (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__A (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__B (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A1 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__B2 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__D (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13669__B1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13309__A1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__D1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__C1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__C1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__B1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__C1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__C1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__B1 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__A1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13315__B1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__A1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__C1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__B1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__S1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__S1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__B1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__C1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__B_N (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__D1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__S0 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14782__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__A1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__A1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__C1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__B1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__C1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__C1 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__A (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__C1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__A (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__C1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13729__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__B1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__C1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13833__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__S0 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13653__S (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__S (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A_N (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__S0 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__S0 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__S0 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__S (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__S0 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__A1 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__A1 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A1 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__S0 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__S0 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S0 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__S0 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12066__A (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__S1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__S1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__B1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__B1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__B1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__B1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__S1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__S1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__S1 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__B1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13740__B1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__A (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14146__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14131__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__C1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__S1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__C1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__C1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A1 (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13930__A1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__B2 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13835__A1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__B2 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__B2 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__C1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__A1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12932__A (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__B2 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A1 (.DIODE(_06425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13659__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__S0 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__A (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__A1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__A_N (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A_N (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__A1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__A1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__A1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__S (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__S (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__C1 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__A (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13835__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__C1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__C1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__A_N (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12510__A (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__S (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__S0 (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A (.DIODE(_06434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13751__A1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__S0 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13657__S1 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__S1 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13622__S1 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__S1 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__S1 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13852__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13718__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__B1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__B1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__S1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__A (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13887__B1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13827__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__S1 (.DIODE(_06438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13614__S (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__S (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13505__S (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A1 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13853__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13758__S (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13629__S (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A1 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A1 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14122__S (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__A (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13932__B2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__B2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13828__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13716__B2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13700__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__B2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__B2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13949__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__B1 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__A1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13716__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__A1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__B2 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__A1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__C1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__C1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__S (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__S (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12166__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A1 (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__A1 (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__S (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13841__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__A (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B2 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__A1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13657__S0 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__S0 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13622__S0 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__S0 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__S0 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13845__S0 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13603__S0 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__S0 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__S0 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__A_N (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13366__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S0 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13851__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13838__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__S (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__S0 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13845__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13603__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__B1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__S1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__A (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13851__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13838__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__C1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__S1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13953__C1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13725__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__A1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13960__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A1 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13371__A (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__S0 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13960__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13639__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__B1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__S1 (.DIODE(_06458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__B1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__B1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__B1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__B1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__C1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__B1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__B1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13936__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13841__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__B1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__B1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__C1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__B1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__B1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__B1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__B1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__C1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__C1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__C1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13569__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__A1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__A1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__B1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__A (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__C1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__B1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__B1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__B2 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__B2 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__C1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A_N (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A1 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13451__A_N (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__A_N (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__S0 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__S (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__S0 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__S0 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__S0 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__B1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__B1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__S1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__S (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__S (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__C1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__S (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__S (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__A (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__A (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__A (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__A (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__C1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__C1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__A (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__A1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__C1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__C1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__A (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13503__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__S0 (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A (.DIODE(_06478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13627__S0 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A1 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__A1 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__S0 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__S (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__S0 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__S0 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__S0 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__B1_N (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__S1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13760__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__B1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__S1 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13535__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13495__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__S (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__S (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__B2 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B2 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__S0 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__A (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__S0 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__A_N (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__A_N (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A_N (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A_N (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__A1 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__S0 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__S (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__S0 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__S0 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13659__S1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__S1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__B1_N (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__B1_N (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__B1_N (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__B1_N (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__S1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12194__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__S1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13488__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__C1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__B1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13663__C1 (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__B1 (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__B1 (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__C1 (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13849__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__B1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__C1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__C1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__C1 (.DIODE(_06497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__B1 (.DIODE(_06497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A (.DIODE(_06497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__A (.DIODE(_06497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A (.DIODE(_06497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__A1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__C1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13729__C1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__B1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__C1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__B1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__C1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__C1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__A1 (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13718__S0 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__A1 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__A_N (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A1 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13361__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A_N (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__S0 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__S0 (.DIODE(_06499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13949__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13935__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__C1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13846__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__B1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__B1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__A (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__A1 (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13703__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__A1 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13538__B_N (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A1 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__S0 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13703__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__B1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__S1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__S0 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__S0 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__S0 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__S0 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__A1 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13950__B_N (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13900__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__S0 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A1 (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__B_N (.DIODE(_06508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13661__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13546__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__B1_N (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__B1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__S1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__A (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__B1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__S1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__B1 (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__S0 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A_N (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A1 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__A (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__S0 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__S0 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__S0 (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__S (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__S (.DIODE(_06514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13953__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__C1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__C1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__B2 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13930__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13840__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13719__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__C1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__C1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13963__A1 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__A1 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__B2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__A1 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A1 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A1 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__S0 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__S0 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__S0 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__S0 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__A1 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__A1 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A1 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__S0 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__B_N (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__S0 (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__S1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__B1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__B1_N (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__A (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12170__A (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__B1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__S1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A2 (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A_N (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13414__A_N (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__A (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12777__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__A (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__S0 (.DIODE(_06527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__B1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13249__B1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12777__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__S1 (.DIODE(_06528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13959__S (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13250__C1 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__C1 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__A (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__S (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13639__S0 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__A (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A1 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__B_N (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__A1 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A1 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13410__A_N (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__S0 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__S0 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__S0 (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__S0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A2 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__B1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__A (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__C1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13827__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13781__A (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__B_N (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__S0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A2 (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__S (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A1 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__S0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__S0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__S0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__S (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__B_N (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__S0 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12913__S0 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__S0 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__S0 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__S0 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12194__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__B_N (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__A (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__S0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13834__S (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13197__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__S (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__S (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S0 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__S (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13932__C1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13849__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13828__B1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13700__C1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__C1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__B2 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__C1 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14139__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14130__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13936__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13757__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__B1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13855__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__C1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__S1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13228__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__S1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__A_N (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__A_N (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A_N (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13416__A_N (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__S0 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__S0 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S0 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__S0 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__S0 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13907__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13844__S (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__S (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__C1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__S (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__S (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__B (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13796__A (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__A (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__S0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A2 (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13963__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13955__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13848__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13727__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__B1 (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13830__C1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__B1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13905__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A1 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__S0 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A1 (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__B_N (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__B1_N (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__B1_N (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__B1_N (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__B1_N (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__S1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__S1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__S1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__S1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__S1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13650__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__B1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__S1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__B1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A0 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A_N (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__A (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A_N (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A_N (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__A_N (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__S0 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__S0 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__S0 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__B1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__C1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__A1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__B1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__C1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__C1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__C1 (.DIODE(_06589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13861__S0 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__S0 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__A1 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__A_N (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A_N (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A_N (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A_N (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__S0 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__S0 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__S0 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13861__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__B1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__S1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A2 (.DIODE(_06595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13955__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13848__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13727__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__B2 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__B2 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__S0 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__S0 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13757__S0 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__S0 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__S (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__A (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S0 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A3 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13769__B1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__C1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__B1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__B2 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13966__B1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13870__B1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__B1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__C1 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A2 (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__C (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__B (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__B (.DIODE(_06609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14230__A (.DIODE(_06609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__B (.DIODE(_06609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14750__A (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__C1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__C1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__B1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__A (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__B1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__B1_N (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__B1_N (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__S1 (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__A (.DIODE(_06614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13751__B1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__B1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__S1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__S1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__S1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__B1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__S1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__C1 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13608__S (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A_N (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__A (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__S0 (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__S0 (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__S (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__S0 (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__S0 (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__S (.DIODE(_06617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__A1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__B1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__B1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__B1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__B1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__B1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__C1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__A (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__C1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__C1 (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13482__C1 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__C1 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__A1 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__A1 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__A1 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13655__A1 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__A (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__A1_N (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__B2 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__A (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A1 (.DIODE(_06624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__A (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__S (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__A1 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__B_N (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__S0 (.DIODE(_06625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13503__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__B1_N (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__S1 (.DIODE(_06627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__B (.DIODE(_06628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__B1 (.DIODE(_06629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13655__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__B1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__B1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__B1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__C1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__A (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__C1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__A (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__B1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13423__C1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__C1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A1 (.DIODE(_06634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A2 (.DIODE(_06635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__B (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__B1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__C1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__B1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__B1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__B1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__C1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__C1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__C1 (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__C1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__C1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__B1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__B1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__B1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__B1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__C1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__B1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__C1 (.DIODE(_06643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13843__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13842__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__A (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__A (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__S0 (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A (.DIODE(_06645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__B1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__B1_N (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__S1 (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__C1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__C1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__S1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__S1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__S1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__S1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__S1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__C1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13654__B2 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__B2 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__C1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A1 (.DIODE(_06650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__A (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__C1 (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__C1 (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__C1 (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__C1 (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__C1 (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A (.DIODE(_06655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__B2 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__S (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A1 (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13661__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13546__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__S0 (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A (.DIODE(_06657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13449__A1 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A1 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A1 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__S0 (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A2 (.DIODE(_06659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13654__C1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__B1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__C1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__C1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__C1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__C1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B1 (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__A (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A (.DIODE(_06660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B (.DIODE(_06661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13509__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__B1 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__B1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13220__B1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__B1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__B1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__C1 (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__A1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13567__A (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__B1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__A (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__A (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__C1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__C1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__C1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__A1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A1 (.DIODE(_06668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__S0 (.DIODE(_06673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__B1 (.DIODE(_06676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__B1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__B1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__C1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__C1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__B2 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__B1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A1 (.DIODE(_06679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__B1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__C1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__C1 (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13375__A (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__C1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A1 (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A1 (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13433__C1 (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__C1 (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__C1 (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__B1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__B1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__B1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__B1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__C1 (.DIODE(_06686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A2 (.DIODE(_06687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__A (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A1 (.DIODE(_06688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A1 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__A1 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__A1 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A1 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__A1 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__S0 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__S0 (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__B1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__B1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__B1_N (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__B1_N (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__B1_N (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__S1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__S1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__B1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__S1 (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__A (.DIODE(_06690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__B1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__S1 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A2 (.DIODE(_06692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__S0 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13785__A (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__S0 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__S0 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13211__A (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A1 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__S0 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__S0 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B_N (.DIODE(_06693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13427__B1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__B1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__B1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__S1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__S1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__S1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__S1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__B1 (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13480__A_N (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A_N (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A_N (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13340__A (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__A1 (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__S0 (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__S (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__S (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__C1 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__B2 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__B2 (.DIODE(_06699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__B1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__B1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__B1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__C1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__C1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__C1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__C1 (.DIODE(_06701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__B1_N (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__B1_N (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__B1_N (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__S1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A0 (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13894__A (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__C1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__B1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__A (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__B1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A1 (.DIODE(_06709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13917__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__S (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__S (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__S0 (.DIODE(_06710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__B1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B1_N (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__B1_N (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__S1 (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A2 (.DIODE(_06712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__B1 (.DIODE(_06713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__B1 (.DIODE(_06716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__S0 (.DIODE(_06717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__B1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__B1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__B1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__S1 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__C1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__C1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__A (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__A (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__C1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__A1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A1 (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__S1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__S1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13449__B1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__B1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__B1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B1_N (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__S1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__S1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__S1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__B1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13517__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__C1 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__B2 (.DIODE(_06728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__B1 (.DIODE(_06729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__S (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13569__A1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13509__A1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__C1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__S (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__S (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__A (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__B1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__B1_N (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__S1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__S1 (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A2 (.DIODE(_06732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__C1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__C1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__A1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__B1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__B1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__B1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__B1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__C1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A1 (.DIODE(_06735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A2 (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13550__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13488__B1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__C1 (.DIODE(_06743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A3 (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A2 (.DIODE(_06746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A2 (.DIODE(_06746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A2 (.DIODE(_06746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__B2 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__A (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__A (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__A2 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A3 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A2 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A2 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__B (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__A2 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__B1 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__B (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A2 (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13573__A (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__C (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A1 (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A1 (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A2 (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A1 (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__B (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A2 (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__B (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A3 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__B (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__A3 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B1 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__C (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A3 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A3 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A1 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A4 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__A2 (.DIODE(_06766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__A0 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__B1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__B1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__B1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__B1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__C1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__D1 (.DIODE(_06769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__B (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__A2 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__B2 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__B1 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__B (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__A2 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__A2 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A2 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__C (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A3 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__A2 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__A2 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A3 (.DIODE(_06781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__B2 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__C (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A2 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__C (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B1 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A2 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14149__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14109__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14067__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__B1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13769__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A1 (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14147__B1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14136__B1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14093__B1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__B1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__A1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__B2 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__A1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__A1 (.DIODE(_06793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A0 (.DIODE(_06794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__S0 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__S0 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__A1 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A_N (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__A_N (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A_N (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__A1 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__A (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__S0 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__S0 (.DIODE(_06795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13812__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__S (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13604__S (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__C1 (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__A1 (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__S (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13427__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__A_N (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__S (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__S0 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__A1 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S0 (.DIODE(_06801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__C1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__C1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__A1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__A1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__A1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__C1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__C1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__C1 (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__S0 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__S0 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__S0 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A1 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A1 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A1 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__A1 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__A1 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__S0 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__S0 (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13627__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__B1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__B1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__S1 (.DIODE(_06811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__B (.DIODE(_06812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__B (.DIODE(_06816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A2 (.DIODE(_06823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__S (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__B2 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__A1 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A1 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A1 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__B2 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__B2 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__A (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A1 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A1 (.DIODE(_06824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A2 (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__A1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__B2 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13327__C1 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__B2 (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A2 (.DIODE(_06834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A2 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__A1 (.DIODE(_06841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__A1 (.DIODE(_06841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__A1 (.DIODE(_06841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13650__S0 (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__S0 (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__A1 (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__A1 (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__A_N (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__A_N (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A_N (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A_N (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__S (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S0 (.DIODE(_06848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A2 (.DIODE(_06849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__B (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__C1 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__B1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13663__A1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__C1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__A1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13550__A1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__C1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__C1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__B1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__C1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A2 (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__S (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__S (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__A1 (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A_N (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__A_N (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__A1 (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__A (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__A1 (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__S0 (.DIODE(_06870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A3 (.DIODE(_06884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13967__B2 (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__A1_N (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__B (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__B1 (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A1 (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B2 (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A3 (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__B (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__A2 (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A2 (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A2_N (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__A1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13284__B1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__C1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__B (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__A (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__B1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__A1 (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A (.DIODE(_06902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__B1 (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__C (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__C (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13285__A (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__B2 (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__B1 (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__B1 (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__B1 (.DIODE(_06910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__B1 (.DIODE(_06916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__B1 (.DIODE(_06916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__B1 (.DIODE(_06916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__A (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__B (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__C1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13779__C1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13585__B1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__B1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__B1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__B1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__C1 (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A1_N (.DIODE(_06918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__B1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__A1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__C (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__A1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__C1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__A1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__C1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__C1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A1 (.DIODE(_06919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__A (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__B1 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13282__A2 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A1 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A1 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__A2 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__A1 (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13674__B1 (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A2 (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A2 (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__B1 (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__A2 (.DIODE(_06923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__B2 (.DIODE(_06938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A2_N (.DIODE(_06938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14115__C1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__C1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__C1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A1 (.DIODE(_06939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__A0 (.DIODE(_06940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__C1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13220__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__A (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__C1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__A1 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__S (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__S (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A1 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A1 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__S (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__S0 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__S0 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__S0 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__S0 (.DIODE(_06946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14071__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__S (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__S (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13855__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__S0 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__A1 (.DIODE(_06951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__A1 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__B2 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__C1 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__B2 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__A (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__A (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__A1 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__B2 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B2 (.DIODE(_06954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__S0 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__S0 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A1 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13263__A (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A_N (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__A1 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A1 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__S (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__S0 (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__B (.DIODE(_06957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__S (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A1 (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13228__A1 (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A1 (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A_N (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A1 (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__S (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__S (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__S (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__S0 (.DIODE(_06959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B (.DIODE(_06961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14149__B1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14067__B1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__C1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__C1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__B1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__B1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13806__C1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__C1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__C1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__C1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__B (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A2 (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13890__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__A1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__A1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12913__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__S1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A2 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__S0 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__S0 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__B_N (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13197__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__S1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__S1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__S0 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__S0 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13852__S0 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__S0 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13651__B_N (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__A_N (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__A_N (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A_N (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__S0 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__S (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A2 (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__S1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13917__S1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__B1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__B1_N (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__B1_N (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__B1_N (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__B1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__S1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__S1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__S1 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A2 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A1_N (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__B1 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14109__B1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__B1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13870__A1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13831__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__A1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13274__C1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__C1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A1 (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A1 (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13900__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__S1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__B1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__S0 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13832__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13752__S (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A1 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A1 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__B_N (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__S0 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S0 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A2 (.DIODE(_07002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13540__S (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__A1 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__S0 (.DIODE(_07008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A2 (.DIODE(_07016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__S0 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13736__S0 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__S0 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__S0 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__A1 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13242__A (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__A (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__S0 (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__A (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__A1 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__S (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__S0 (.DIODE(_07022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A2 (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__B1 (.DIODE(_07037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A3 (.DIODE(_07038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A2 (.DIODE(_07062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A2 (.DIODE(_07062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A2 (.DIODE(_07062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A0 (.DIODE(_07063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A1 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__A (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__A1 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__B2 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__A1 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__B2 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__B2 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__B2 (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A (.DIODE(_07066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13890__S0 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__A1 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__B_N (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A1 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A1 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__B_N (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__S0 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__S0 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__S0 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__B1 (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__B1 (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__B1 (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__S (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B1 (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__C1 (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A (.DIODE(_07070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__B1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13908__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A1 (.DIODE(_07071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__B1_N (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__B1_N (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__B1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__S1 (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A (.DIODE(_07072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13905__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__S1 (.DIODE(_07073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A1 (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14125__S0 (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__S0 (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__S0 (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14015__S0 (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__A (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13910__S (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__S (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__S (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__S (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A1 (.DIODE(_07079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__B (.DIODE(_07083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__C1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__C1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__A1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__A (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__C1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__B1 (.DIODE(_07085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__B (.DIODE(_07087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__B1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__B1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__B1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__B1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__C1 (.DIODE(_07094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A2 (.DIODE(_07095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__S (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A1 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__A1 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__B2 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__B2 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__A (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A1 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A1 (.DIODE(_07096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__S0 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__A1 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13856__B_N (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13740__A1 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13739__B_N (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__A1 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A1 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__S0 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__S0 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S0 (.DIODE(_07097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__S1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__B1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__B1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__B1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__B1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__B1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__S1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__S1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__S1 (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A (.DIODE(_07098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__A (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S1 (.DIODE(_07099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A2 (.DIODE(_07100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__B2 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__C1 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__B2 (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__A1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13908__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__C1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A2 (.DIODE(_07110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13843__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13842__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__B1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__B1_N (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__S1 (.DIODE(_07111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A2 (.DIODE(_07114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__B1 (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__B1 (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__B1 (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A1 (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A2 (.DIODE(_07126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__A (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__B1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__C1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__A1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__C1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__B1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A1 (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A2 (.DIODE(_07137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A2 (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B2 (.DIODE(_07158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__B1 (.DIODE(_07159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A3 (.DIODE(_07160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__S (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13883__S0 (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__S (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A1 (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__S (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__B (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__S (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__S0 (.DIODE(_07164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__B1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__C1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14006__B1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13830__A1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A1 (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__A1 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14115__B2 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__B2 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14040__S (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__S (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__A1 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__B2 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__A1 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A1 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A1 (.DIODE(_07203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14144__S (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14110__A (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14095__A1 (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14094__B_N (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__S (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13981__A (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__S0 (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__S0 (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__S0 (.DIODE(_07204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14143__B1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14063__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14052__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14015__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__A (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__A (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12945__A (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__S1 (.DIODE(_07205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14145__B2 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14113__A1 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__B2 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__A1 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__B2 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__A1 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__B2 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__A1 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13814__A (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A1 (.DIODE(_07207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__S1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14125__S1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14095__B1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__S1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__S1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__A (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__B1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__B1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__B1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__B1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__C1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__C1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__C1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__C1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__C1 (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__A (.DIODE(_07219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14132__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14126__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__A (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__B1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__A1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__C1 (.DIODE(_07220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13245__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A1 (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13929__S (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__A1 (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13249__A1 (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__A1 (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__S (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__S (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__S (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__S (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__A (.DIODE(_07227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__B1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A2 (.DIODE(_07235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__B (.DIODE(_07236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A2 (.DIODE(_07238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__B (.DIODE(_07240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__B (.DIODE(_07245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A2 (.DIODE(_07248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A3 (.DIODE(_07253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14106__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14080__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13833__C1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__S1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__C1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A1 (.DIODE(_07257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13760__S0 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__S0 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__S0 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A1 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A1 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A1 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A_N (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A_N (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__S0 (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__S (.DIODE(_07263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A2 (.DIODE(_07275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__B1 (.DIODE(_07280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__A2_N (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__B (.DIODE(_07289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__B1 (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__B1 (.DIODE(_07311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A3 (.DIODE(_07312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A3 (.DIODE(_07312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A3 (.DIODE(_07312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B (.DIODE(_07312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__A1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14172__S0 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14161__A1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14160__B1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__S1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__S1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__A1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__B1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__A1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A1 (.DIODE(_07322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__B1 (.DIODE(_07337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A2 (.DIODE(_07338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A2 (.DIODE(_07339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A2 (.DIODE(_07350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__C1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14100__C1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__B1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__B1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A1 (.DIODE(_07354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14105__A (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__C1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13793__B1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A1 (.DIODE(_07355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A0 (.DIODE(_07366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13784__A (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__A (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__A1 (.DIODE(_07376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A1 (.DIODE(_07376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A2 (.DIODE(_07384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13797__A (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13736__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__B1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__S1 (.DIODE(_07391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A2 (.DIODE(_07397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A1 (.DIODE(_07403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A2 (.DIODE(_07408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__B2 (.DIODE(_07416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A3 (.DIODE(_07418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_i_A (.DIODE(clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A1 (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A (.DIODE(\fifo0.fifo_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A1 (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A (.DIODE(\fifo0.fifo_data[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A1 (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__A (.DIODE(\fifo0.fifo_data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11418__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A1 (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__A (.DIODE(\fifo0.fifo_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__A1 (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A (.DIODE(\fifo0.fifo_data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A1 (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A (.DIODE(\fifo0.fifo_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A1 (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__A (.DIODE(\fifo0.fifo_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A1 (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A (.DIODE(\fifo0.fifo_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A1 (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A (.DIODE(\fifo0.fifo_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A1 (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A (.DIODE(\fifo0.fifo_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A1 (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A (.DIODE(\fifo0.fifo_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__A1 (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A (.DIODE(\fifo0.fifo_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__A2 (.DIODE(\fifo0.fifo_store[106][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A0 (.DIODE(\fifo0.fifo_store[106][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__A1 (.DIODE(\fifo0.fifo_store[45][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A0 (.DIODE(\fifo0.fifo_store[45][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__A1 (.DIODE(\fifo0.fifo_store[45][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A0 (.DIODE(\fifo0.fifo_store[45][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13657__A1 (.DIODE(\fifo0.fifo_store[49][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A0 (.DIODE(\fifo0.fifo_store[49][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(fifo_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(fifo_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(fifo_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(fifo_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(fifo_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(fifo_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(fifo_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(fifo_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(fifo_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(fifo_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(fifo_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(fifo_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(fifo_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(fifo_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(fifo_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(fifo_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(fifo_rdy_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(mode_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(osr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(osr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(rst_n_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(tst_fifo_loop_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(tst_sinegen_en_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(tst_sinegen_step_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(tst_sinegen_step_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(tst_sinegen_step_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(tst_sinegen_step_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(tst_sinegen_step_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(tst_sinegen_step_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(volume_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(volume_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(volume_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(volume_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__C1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__C1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__14753__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__14759__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__14761__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__14760__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__14773__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__14782__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__C1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__13878__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__C1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__14173__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__13973__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__D (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__D (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_i_A (.DIODE(clknet_1_0_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_i_A (.DIODE(clknet_1_0_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_i_A (.DIODE(clknet_1_1_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_i_A (.DIODE(clknet_1_1_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_i_A (.DIODE(clknet_2_0_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_i_A (.DIODE(clknet_2_0_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_i_A (.DIODE(clknet_2_1_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_i_A (.DIODE(clknet_2_1_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_i_A (.DIODE(clknet_2_2_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_i_A (.DIODE(clknet_2_2_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_i_A (.DIODE(clknet_2_3_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_i_A (.DIODE(clknet_2_3_1_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_i_A (.DIODE(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_i_A (.DIODE(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_i_A (.DIODE(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_i_A (.DIODE(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_i_A (.DIODE(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_i_A (.DIODE(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_i_A (.DIODE(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_i_A (.DIODE(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_i_A (.DIODE(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_i_A (.DIODE(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_i_A (.DIODE(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_i_A (.DIODE(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_i_A (.DIODE(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_i_A (.DIODE(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_i_A (.DIODE(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_i_A (.DIODE(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_1_0_clk_i_A (.DIODE(clknet_4_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_0_0_clk_i_A (.DIODE(clknet_4_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_3_0_clk_i_A (.DIODE(clknet_4_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_2_0_clk_i_A (.DIODE(clknet_4_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_5_0_clk_i_A (.DIODE(clknet_4_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_4_0_clk_i_A (.DIODE(clknet_4_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_7_0_clk_i_A (.DIODE(clknet_4_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_6_0_clk_i_A (.DIODE(clknet_4_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_9_0_clk_i_A (.DIODE(clknet_4_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_8_0_clk_i_A (.DIODE(clknet_4_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_11_0_clk_i_A (.DIODE(clknet_4_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_10_0_clk_i_A (.DIODE(clknet_4_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_13_0_clk_i_A (.DIODE(clknet_4_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_12_0_clk_i_A (.DIODE(clknet_4_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_15_0_clk_i_A (.DIODE(clknet_4_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_14_0_clk_i_A (.DIODE(clknet_4_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_17_0_clk_i_A (.DIODE(clknet_4_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_16_0_clk_i_A (.DIODE(clknet_4_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_19_0_clk_i_A (.DIODE(clknet_4_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_18_0_clk_i_A (.DIODE(clknet_4_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_21_0_clk_i_A (.DIODE(clknet_4_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_20_0_clk_i_A (.DIODE(clknet_4_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_23_0_clk_i_A (.DIODE(clknet_4_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_22_0_clk_i_A (.DIODE(clknet_4_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_25_0_clk_i_A (.DIODE(clknet_4_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_24_0_clk_i_A (.DIODE(clknet_4_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_27_0_clk_i_A (.DIODE(clknet_4_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_26_0_clk_i_A (.DIODE(clknet_4_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_29_0_clk_i_A (.DIODE(clknet_4_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_28_0_clk_i_A (.DIODE(clknet_4_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_31_0_clk_i_A (.DIODE(clknet_4_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_30_0_clk_i_A (.DIODE(clknet_4_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_341_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_340_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_339_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_338_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_337_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_i_A (.DIODE(clknet_5_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_343_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_342_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_336_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_335_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__CLK (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_333_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_329_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_i_A (.DIODE(clknet_5_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_i_A (.DIODE(clknet_5_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_i_A (.DIODE(clknet_5_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_332_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_331_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_330_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_328_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_327_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_326_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_315_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_314_clk_i_A (.DIODE(clknet_5_4_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_325_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_324_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_323_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_322_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_321_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_320_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_319_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_318_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_317_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_316_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_308_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_307_clk_i_A (.DIODE(clknet_5_5_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_313_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_312_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_311_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_i_A (.DIODE(clknet_5_6_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_310_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_309_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_306_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_305_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_304_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_303_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_302_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_i_A (.DIODE(clknet_5_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_i_A (.DIODE(clknet_5_8_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_i_A (.DIODE(clknet_5_9_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_i_A (.DIODE(clknet_5_10_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_i_A (.DIODE(clknet_5_11_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_i_A (.DIODE(clknet_5_12_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_i_A (.DIODE(clknet_5_13_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_i_A (.DIODE(clknet_5_14_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_i_A (.DIODE(clknet_5_15_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_285_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_284_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_283_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_282_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_281_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_280_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_279_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_278_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_277_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__CLK (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_275_clk_i_A (.DIODE(clknet_5_16_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_289_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_287_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_286_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_274_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_273_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_272_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_271_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_270_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_269_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_268_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_267_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_266_clk_i_A (.DIODE(clknet_5_17_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_301_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_300_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_299_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_298_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_297_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_296_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_295_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_220_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_219_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_218_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_217_clk_i_A (.DIODE(clknet_5_18_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_294_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_293_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_292_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_291_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_290_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_288_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_225_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_221_clk_i_A (.DIODE(clknet_5_19_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_265_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_264_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_263_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_262_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_261_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_260_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_259_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_253_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_251_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_250_clk_i_A (.DIODE(clknet_5_20_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_258_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_257_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_256_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_255_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_254_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_252_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_249_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_246_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_245_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_244_clk_i_A (.DIODE(clknet_5_21_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_234_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_233_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_232_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_231_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_230_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_229_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_228_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_227_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_226_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_224_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_223_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_222_clk_i_A (.DIODE(clknet_5_22_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_248_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_247_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_243_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_242_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_241_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_240_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_239_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_238_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_237_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_236_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_235_clk_i_A (.DIODE(clknet_5_23_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_216_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_215_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_214_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_213_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_i_A (.DIODE(clknet_5_24_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_212_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_211_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_210_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_208_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_207_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_206_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_205_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_i_A (.DIODE(clknet_5_25_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_i_A (.DIODE(clknet_5_26_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_i_A (.DIODE(clknet_5_27_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_209_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_203_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_202_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_201_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_200_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_199_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_198_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_197_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_196_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_195_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_194_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_193_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_i_A (.DIODE(clknet_5_28_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_192_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_191_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_189_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_i_A (.DIODE(clknet_5_29_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_204_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_i_A (.DIODE(clknet_5_30_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_i_A (.DIODE(clknet_5_31_0_clk_i));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1311 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1334 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1318 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1423 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1282 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1334 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1362 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1327 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1422 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1288 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1395 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1290 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1309 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1334 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1280 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1393 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1396 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1260 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1307 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1404 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1375 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1312 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1380 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1387 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1396 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1372 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1422 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1417 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1292 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1346 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1306 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1362 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1404 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1280 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1288 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1419 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1368 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1293 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1380 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1376 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1422 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1362 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1375 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1388 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1376 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1419 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1396 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1386 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1392 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1384 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1306 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1334 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1330 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1360 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1316 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1339 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1347 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1277 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1344 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1388 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1417 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1339 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1380 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1264 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1324 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1386 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1334 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1346 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1291 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1334 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1337 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1284 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1413 ();
endmodule

